** sch_path: /home/designer/shared/Workshop-CANELOS24/xschem/TB_hvNMOS_charact.sch
**.subckt TB_hvNMOS_charact
XM1 net1 Vg GND GND sg13_hv_nmos w={w_M1} l={l_M1} ng=1 m={mult_M1}
Vgs Vg GND 3.3
Vds Vd GND 3
VdM1 Vd net1 0
.save i(vdm1)
XM2 net2 Vg GND GND sg13_hv_nmos w={w_M2} l={l_M2} ng=1 m={mult_M2}
VdM2 Vd net2 0
.save i(vdm2)
XM3 net3 Vg GND GND sg13_hv_nmos w={w_M3} l={l_M3} ng=1 m={mult_M3}
VdM3 Vd net3 0
.save i(vdm3)
**** begin user architecture code


.param temp=27
.param mult_M1 = 1200
.param w_M1 =10u
.param l_M1 =0.22u

.param mult_M2 = 1200
.param w_M2 =10u
.param l_M2 =0.25u

.param mult_M3 = 1200
.param w_M3 =10u
.param l_M3 =0.35u

.save all
* + @M.XM1.m1[id]
+ @n.xm1.nsg13_hv_nmos[vth]
+ @n.xm1.nsg13_hv_nmos[gds]
+ @n.xm2.nsg13_hv_nmos[vth]
+ @n.xm2.nsg13_hv_nmos[gds]
+ @n.xm3.nsg13_hv_nmos[vth]
+ @n.xm3.nsg13_hv_nmos[gds]
+ @n.xm1.nsg13_hv_nmos[ad]

.control
*dc Vds 0 3 0.01 Vgs 0.5 3 0.5
dc Vds 0 3 0.01
*dc Vds 0 0.5 0.01
*dc Vds 0 0.5 0.01 temp 0 27 1
write dc_hv_nmos.raw
let G_M1 = @n.xm1.nsg13_hv_nmos[gds]
let G_M2 = @n.xm2.nsg13_hv_nmos[gds]
let G_M3 = @n.xm3.nsg13_hv_nmos[gds]
let Ron_M1 = 1/G_M1
let Ron_M2 = 1/G_M2
let Ron_M3 = 1/G_M3
let Vds = v(Vd)

let Vth_M1 = @n.xm1.nsg13_hv_nmos[vth]
let Id_M1 = i(VdM1)
plot i(VdM1) i(VdM2) i(VdM3) vs Vds
plot Ron_M1 Ron_M2 Ron_M3 vs Vds
*plot Id_M1
*plot Vth_M1 Vth_M1*2
*print @n.xm1.nsg13_hv_nmos[vth] @n.xm2.nsg13_hv_nmos[vth] Vth_M1
*print @n.xm2.nsg13_hv_nmos[vth]
write test_nmos.raw




.endc



.lib cornerMOShv.lib mos_tt

**** end user architecture code
**.ends
.GLOBAL GND
.end
