module tb_grid;

    // Inputs
    reg [7:0] din;
    reg [7:0] sign;  // Single 8-bit vector
    reg [7:0] win0, win1, win2, win3, win4, win5, win6, win7;  // Individual inputs for win
    reg [7:0] bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7;  // Individual inputs for bias
    reg trig;
    reg clk;
    reg rst;

    // Outputs
    wire [7:0] dout0, dout1, dout2, dout3, dout4, dout5, dout6, dout7;  // Individual outputs

    // Instantiate the Unit Under Test (UUT)
    grid uut (
        .din(din),
        .sign(sign),  // Single sign input
        .win0(win0), .win1(win1), .win2(win2), .win3(win3),
        .win4(win4), .win5(win5), .win6(win6), .win7(win7),
        .bias0(bias0), .bias1(bias1), .bias2(bias2), .bias3(bias3),
        .bias4(bias4), .bias5(bias5), .bias6(bias6), .bias7(bias7),
        .dout0(dout0), .dout1(dout1), .dout2(dout2), .dout3(dout3),
        .dout4(dout4), .dout5(dout5), .dout6(dout6), .dout7(dout7),
        .trig(trig),
        .clk(clk),
        .rst(rst)
    );

    // Clock generation
    initial begin
        clk = 0;
        forever #5 clk = ~clk;  // Clock with a period of 10 time units
    end

    // Test stimulus
    initial begin
        // Open VCD file for waveform viewing
        $dumpfile("results/tb_grid.vcd");
        $dumpvars(0, tb_grid);

        // Monitor output
        $monitor("Time: %0d | din: %d | trig: %b | rst: %b | dout0: %d | dout1: %d | dout2: %d | dout3: %d | dout4: %d | dout5: %d | dout6: %d | dout7: %d",
                 $time, din, trig, rst, dout0, dout1, dout2, dout3, dout4, dout5, dout6, dout7);

        // Initialize inputs
        rst = 1;
        din = 8'd0;
        trig = 0;

        // Initialize sign, win, and bias
        sign = 8'b00000000;

        win0 = 8'd0; win1 = 8'd0; win2 = 8'd0; win3 = 8'd0;
        win4 = 8'd0; win5 = 8'd0; win6 = 8'd0; win7 = 8'd0;

        bias0 = 8'd0; bias1 = 8'd0; bias2 = 8'd0; bias3 = 8'd0;
        bias4 = 8'd0; bias5 = 8'd0; bias6 = 8'd0; bias7 = 8'd0;

        #20 rst = 0;  // Release reset

        // Operation 1: 
        // x=32, 
        // s=[-1.  1. -1.  1.  1. -1.  1. -1.],
        // w=[ 7  9  3  0 11  7  6  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-224.  288.  -96.    0.  352. -224.  192.  -64.], 
        // Q{mac}=[0 0 0 0 0 0 0 0]

        sign=8'b01011010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00001001, 8'b00000011, 8'b00000000, 8'b00001011, 8'b00000111, 8'b00000110, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00100000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 2: 
        // x=-4, 
        // s=[ 1.  1. -1.  1.  1. -1. -1.  1.],
        // w=[17 45 34  2 23 32 17  6],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-292.  108.   40.   -8.  260.  -96.  260.  -88.], 
        // Q{mac}=[0 0 0 0 0 0 0 0]

        sign=8'b11011001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00010001, 8'b00101101, 8'b00100010, 8'b00000010, 8'b00010111, 8'b00100000, 8'b00010001, 8'b00000110};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11111100;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 3: 
        // x=-3, 
        // s=[-1. -1. -1.  1.  1. -1.  1.  1.],
        // w=[ 2  1 11  6 25 19  3  7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-286.  111.   73.  -26.  185.  -39.  251. -109.], 
        // Q{mac}=[0 0 0 0 0 0 0 0]

        sign=8'b00011011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00000001, 8'b00001011, 8'b00000110, 8'b00011001, 8'b00010011, 8'b00000011, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11111101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 4: 
        // x=-121, 
        // s=[ 1.  1. -1. -1. -1.  1.  1.  1.],
        // w=[ 4 12 14 19  7 20 13  9],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -770. -1341.  1767.  2273.  1032. -2459. -1322. -1198.], 
        // Q{mac}=[0 0 1 2 1 0 0 0]

        sign=8'b11000111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000100, 8'b00001100, 8'b00001110, 8'b00010011, 8'b00000111, 8'b00010100, 8'b00001101, 8'b00001001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000111;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 5: 
        // x=-118, 
        // s=[-1. -1.  1.  1.  1.  1.  1.  1.],
        // w=[15 11  9  8 12 11  4  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 1000.   -43.   705.  1329.  -384. -3757. -1794. -1552.], 
        // Q{mac}=[0 0 0 1 0 0 0 0]

        sign=8'b00111111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001111, 8'b00001011, 8'b00001001, 8'b00001000, 8'b00001100, 8'b00001011, 8'b00000100, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 6: 
        // x=-86, 
        // s=[-1. -1.  1.  1.  1.  1.  1.  1.],
        // w=[3 2 9 4 6 6 5 5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 1258.   129.   -69.   985.  -900. -4273. -2224. -1982.], 
        // Q{mac}=[1 0 0 0 0 0 0 0]

        sign=8'b00111111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00000010, 8'b00001001, 8'b00000100, 8'b00000110, 8'b00000110, 8'b00000101, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10101010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 7: 
        // x=-122, 
        // s=[ 1.  1. -1. -1.  1.  1. -1.  1.],
        // w=[ 7 12  7 21 10 15  1  1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  404. -1335.   785.  3547. -2120. -6103. -2102. -2104.], 
        // Q{mac}=[0 0 0 3 0 0 0 0]

        sign=8'b11001101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00001100, 8'b00000111, 8'b00010101, 8'b00001010, 8'b00001111, 8'b00000001, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 8: 
        // x=-119, 
        // s=[-1. -1.  1.  1.  1.  1. -1.  1.],
        // w=[17 11  7  0  5  5  3  9],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 2427.   -26.   -48.  3547. -2715. -6698. -1745. -3175.], 
        // Q{mac}=[2 0 0 3 0 0 0 0]

        sign=8'b00111101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00010001, 8'b00001011, 8'b00000111, 8'b00000000, 8'b00000101, 8'b00000101, 8'b00000011, 8'b00001001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 9: 
        // x=-87, 
        // s=[-1. -1.  1. -1. -1.  1.  1.  1.],
        // w=[15 12  0  2  5  8  4  7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 3732.  1018.   -48.  3721. -2280. -7394. -2093. -3784.], 
        // Q{mac}=[3 0 0 3 0 0 0 0]

        sign=8'b00100111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001111, 8'b00001100, 8'b00000000, 8'b00000010, 8'b00000101, 8'b00001000, 8'b00000100, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10101001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 10: 
        // x=-115, 
        // s=[ 1.  1. -1. -1.  1.  1.  1.  1.],
        // w=[ 2 18 24 30 10  9 17  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 3502. -1052.  2712.  7171. -3430. -8429. -4048. -4359.], 
        // Q{mac}=[3 0 2 7 0 0 0 0]

        sign=8'b11001111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00010010, 8'b00011000, 8'b00011110, 8'b00001010, 8'b00001001, 8'b00010001, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 11: 
        // x=-72, 
        // s=[-1. -1.  1. -1. -1.  1.  1.  1.],
        // w=[ 1  7 15  3 10 20  1  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 3574.  -548.  1632.  7387. -2710. -9869. -4120. -4575.], 
        // Q{mac}=[3 0 1 7 0 0 0 0]

        sign=8'b00100111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00000111, 8'b00001111, 8'b00000011, 8'b00001010, 8'b00010100, 8'b00000001, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10111000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 12: 
        // x=-60, 
        // s=[-1. -1. -1.  1. -1.  1.  1.  1.],
        // w=[12  1  2  3  9 11  3  8],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  4294.   -488.   1752.   7207.  -2170. -10529.  -4300.  -5055.], 
        // Q{mac}=[4 0 1 7 0 0 0 0]

        sign=8'b00010111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001100, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00001001, 8'b00001011, 8'b00000011, 8'b00001000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11000100;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 13: 
        // x=90, 
        // s=[ 1.  1. -1.  1.  1. -1. -1. -1.],
        // w=[ 7  5  4 11 19 17 11  7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  4924.    -38.   1392.   8197.   -460. -12059.  -5290.  -5685.], 
        // Q{mac}=[4 0 1 8 0 0 0 0]

        sign=8'b11011000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00000101, 8'b00000100, 8'b00001011, 8'b00010011, 8'b00010001, 8'b00001011, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b01011010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 14: 
        // x=80, 
        // s=[ 1.  1.  1.  1. -1. -1.  1. -1.],
        // w=[12  7  5  8 12 15  0 11],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  5884.    522.   1792.   8837.  -1420. -13259.  -5290.  -6565.], 
        // Q{mac}=[5 0 1 8 0 0 0 0]

        sign=8'b11110010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001100, 8'b00000111, 8'b00000101, 8'b00001000, 8'b00001100, 8'b00001111, 8'b00000000, 8'b00001011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b01010000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 15: 
        // x=100, 
        // s=[ 1. -1.  1. -1. -1. -1. -1.  1.],
        // w=[0 6 7 3 9 3 1 1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  5884.    -78.   2492.   8537.  -2320. -13559.  -5390.  -6465.], 
        // Q{mac}=[5 0 2 8 0 0 0 0]

        sign=8'b10100001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000000, 8'b00000110, 8'b00000111, 8'b00000011, 8'b00001001, 8'b00000011, 8'b00000001, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b01100100;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 16: 
        // x=-113, 
        // s=[-1.  1. -1. -1.  1.  1.  1. -1.],
        // w=[ 9 10  7 11  6 17  6  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  6901.  -1208.   3283.   9780.  -2998. -15480.  -6068.  -5900.], 
        // Q{mac}=[6 0 3 9 0 0 0 0]

        sign=8'b01001110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001001, 8'b00001010, 8'b00000111, 8'b00001011, 8'b00000110, 8'b00010001, 8'b00000110, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001111;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 17: 
        // x=-128, 
        // s=[ 1.  1. -1. -1.  1.  1.  1.  1.],
        // w=[ 0 10 17  8  4  1  4  7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  6901.  -2488.   5459.  10804.  -3510. -15608.  -6580.  -6796.], 
        // Q{mac}=[ 6  0  5 10  0  0  0  0]

        sign=8'b11001111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000000, 8'b00001010, 8'b00010001, 8'b00001000, 8'b00000100, 8'b00000001, 8'b00000100, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 18: 
        // x=-128, 
        // s=[ 1. -1.  1.  1.  1.  1. -1.  1.],
        // w=[ 0 10  2  1  2  1  2  0],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  6901.  -1208.   5203.  10676.  -3766. -15736.  -6324.  -6796.], 
        // Q{mac}=[ 6  0  5 10  0  0  0  0]

        sign=8'b10111101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000000, 8'b00001010, 8'b00000010, 8'b00000001, 8'b00000010, 8'b00000001, 8'b00000010, 8'b00000000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 19: 
        // x=-120, 
        // s=[-1.  1. -1.  1. -1.  1.  1. -1.],
        // w=[2 5 8 0 3 1 4 1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  7141.  -1808.   6163.  10676.  -3406. -15856.  -6804.  -6676.], 
        // Q{mac}=[ 6  0  6 10  0  0  0  0]

        sign=8'b01010110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00000101, 8'b00001000, 8'b00000000, 8'b00000011, 8'b00000001, 8'b00000100, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 20: 
        // x=-125, 
        // s=[ 1.  1.  1. -1.  1.  1. -1. -1.],
        // w=[ 4  5  1 10  7  5  2  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  6641.  -2433.   6038.  11926.  -4281. -16481.  -6554.  -6051.], 
        // Q{mac}=[ 6  0  5 11  0  0  0  0]

        sign=8'b11101100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000100, 8'b00000101, 8'b00000001, 8'b00001010, 8'b00000111, 8'b00000101, 8'b00000010, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000011;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 21: 
        // x=-122, 
        // s=[-1. -1.  1. -1. -1.  1. -1.  1.],
        // w=[ 3  4  8  2 15  9  6 10],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  7007.  -1945.   5062.  12170.  -2451. -17579.  -5822.  -7271.], 
        // Q{mac}=[ 6  0  4 11  0  0  0  0]

        sign=8'b00100101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00000100, 8'b00001000, 8'b00000010, 8'b00001111, 8'b00001001, 8'b00000110, 8'b00001010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 22: 
        // x=-107, 
        // s=[ 1. -1.  1. -1. -1.  1.  1.  1.],
        // w=[ 0  1  6  1 10  4  5  0],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  7007.  -1838.   4420.  12277.  -1381. -18007.  -6357.  -7271.], 
        // Q{mac}=[ 6  0  4 11  0  0  0  0]

        sign=8'b10100111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000000, 8'b00000001, 8'b00000110, 8'b00000001, 8'b00001010, 8'b00000100, 8'b00000101, 8'b00000000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10010101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 23: 
        // x=-22, 
        // s=[-1. -1.  1.  1. -1.  1.  1.  1.],
        // w=[ 8 25 15 19  1  1  1  1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  7183.  -1288.   4090.  11859.  -1359. -18029.  -6379.  -7293.], 
        // Q{mac}=[ 7  0  3 11  0  0  0  0]

        sign=8'b00110111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001000, 8'b00011001, 8'b00001111, 8'b00010011, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11101010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 24: 
        // x=-49, 
        // s=[ 1.  1. -1. -1.  1. -1. -1.  1.],
        // w=[10 24 11  7 34  4  3  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  6693.  -2464.   4629.  12202.  -3025. -17833.  -6232.  -7538.], 
        // Q{mac}=[ 6  0  4 11  0  0  0  0]

        sign=8'b11001001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001010, 8'b00011000, 8'b00001011, 8'b00000111, 8'b00100010, 8'b00000100, 8'b00000011, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11001111;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 25: 
        // x=30, 
        // s=[ 1.  1. -1. -1.  1. -1. -1.  1.],
        // w=[10 28 27  8 44 30 10  4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  6993.  -1624.   3819.  11962.  -1705. -18733.  -6532.  -7418.], 
        // Q{mac}=[ 6  0  3 11  0  0  0  0]

        sign=8'b11001001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001010, 8'b00011100, 8'b00011011, 8'b00001000, 8'b00101100, 8'b00011110, 8'b00001010, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00011110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 26: 
        // x=65, 
        // s=[ 1. -1. -1.  1.  1. -1.  1.  1.],
        // w=[ 1  6 14  7  2  8 11  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  7058.  -2014.   2909.  12417.  -1575. -19253.  -5817.  -7223.], 
        // Q{mac}=[ 6  0  2 12  0  0  0  0]

        sign=8'b10011011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00000110, 8'b00001110, 8'b00000111, 8'b00000010, 8'b00001000, 8'b00001011, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b01000001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 27: 
        // x=-63, 
        // s=[-1. -1.  1.  1.  1.  1. -1. -1.],
        // w=[11 22 14  4  0  5 16  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  7751.   -628.   2027.  12165.  -1575. -19568.  -4809.  -7034.], 
        // Q{mac}=[ 7  0  1 11  0  0  0  0]

        sign=8'b00111100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001011, 8'b00010110, 8'b00001110, 8'b00000100, 8'b00000000, 8'b00000101, 8'b00010000, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11000001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 28: 
        // x=60, 
        // s=[-1.  1.  1.  1.  1.  1. -1.  1.],
        // w=[ 7  2 11  6  3  3 15  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  7331.   -508.   2687.  12525.  -1395. -19388.  -5709.  -6914.], 
        // Q{mac}=[ 7  0  2 12  0  0  0  0]

        sign=8'b01111101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00000010, 8'b00001011, 8'b00000110, 8'b00000011, 8'b00000011, 8'b00001111, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00111100;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 29: 
        // x=-7, 
        // s=[ 1.  1. -1. -1.  1. -1.  1. -1.],
        // w=[28 35 42 30 16 17  7  4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  7135.   -753.   2981.  12735.  -1507. -19269.  -5758.  -6886.], 
        // Q{mac}=[ 6  0  2 12  0  0  0  0]

        sign=8'b11001010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00011100, 8'b00100011, 8'b00101010, 8'b00011110, 8'b00010000, 8'b00010001, 8'b00000111, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11111001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 30: 
        // x=26, 
        // s=[-1.  1. -1. -1.  1. -1.  1. -1.],
        // w=[ 3  9 11 11  7 19  5 10],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  7057.   -519.   2695.  12449.  -1325. -19763.  -5628.  -7146.], 
        // Q{mac}=[ 6  0  2 12  0  0  0  0]

        sign=8'b01001010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00001001, 8'b00001011, 8'b00001011, 8'b00000111, 8'b00010011, 8'b00000101, 8'b00001010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00011010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 31: 
        // x=-18, 
        // s=[-1.  1.  1.  1. -1.  1. -1.  1.],
        // w=[ 1  7  1 12  6 19  7  9],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  7075.   -645.   2677.  12233.  -1217. -20105.  -5502.  -7308.], 
        // Q{mac}=[ 6  0  2 11  0  0  0  0]

        sign=8'b01110101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00000111, 8'b00000001, 8'b00001100, 8'b00000110, 8'b00010011, 8'b00000111, 8'b00001001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11101110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 32: 
        // x=16, 
        // s=[-1. -1. -1. -1.  1. -1.  1. -1.],
        // w=[ 2  5  6  4 10  7  4 14],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  7043.   -725.   2581.  12169.  -1057. -20217.  -5438.  -7532.], 
        // Q{mac}=[ 6  0  2 11  0  0  0  0]

        sign=8'b00001010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00000101, 8'b00000110, 8'b00000100, 8'b00001010, 8'b00000111, 8'b00000100, 8'b00001110};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00010000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 33: 
        // x=-3, 
        // s=[ 1.  1. -1. -1.  1. -1. -1.  1.],
        // w=[25 42  1 23 16  8 36  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  6968.   -851.   2584.  12238.  -1105. -20193.  -5330.  -7538.], 
        // Q{mac}=[ 6  0  2 11  0  0  0  0]

        sign=8'b11001001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00011001, 8'b00101010, 8'b00000001, 8'b00010111, 8'b00010000, 8'b00001000, 8'b00100100, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11111101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 34: 
        // x=-15, 
        // s=[-1. -1. -1.  1.  1. -1.  1.  1.],
        // w=[ 2 10  8  2  7 23 17  6],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  6998.   -701.   2704.  12208.  -1210. -19848.  -5585.  -7628.], 
        // Q{mac}=[ 6  0  2 11  0  0  0  0]

        sign=8'b00011011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00001010, 8'b00001000, 8'b00000010, 8'b00000111, 8'b00010111, 8'b00010001, 8'b00000110};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11110001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 35: 
        // x=8, 
        // s=[-1.  1. -1.  1.  1. -1.  1.  1.],
        // w=[ 3  3  2  3 17  7  1  4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  6974.   -677.   2688.  12232.  -1074. -19904.  -5577.  -7596.], 
        // Q{mac}=[ 6  0  2 11  0  0  0  0]

        sign=8'b01011011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00000011, 8'b00000010, 8'b00000011, 8'b00010001, 8'b00000111, 8'b00000001, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00001000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 36: 
        // x=-23, 
        // s=[ 1.  1.  1. -1.  1.  1.  1.  1.],
        // w=[ 8 11  0  6  0 18  0  4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  6790.   -930.   2688.  12370.  -1074. -20318.  -5577.  -7688.], 
        // Q{mac}=[ 6  0  2 12  0  0  0  0]

        sign=8'b11101111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001000, 8'b00001011, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00010010, 8'b00000000, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11101001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 37: 
        // x=4, 
        // s=[ 1.  1.  1. -1. -1.  1. -1.  1.],
        // w=[36  8 28  1 30 23 31  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  6934.   -898.   2800.  12366.  -1194. -20226.  -5701.  -7680.], 
        // Q{mac}=[ 6  0  2 12  0  0  0  0]

        sign=8'b11100101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00100100, 8'b00001000, 8'b00011100, 8'b00000001, 8'b00011110, 8'b00010111, 8'b00011111, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00000100;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 38: 
        // x=9, 
        // s=[-1. -1.  1.  1. -1. -1. -1. -1.],
        // w=[ 9 14 26 66  7 27 47  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  6853.  -1024.   3034.  12960.  -1257. -20469.  -6124.  -7725.], 
        // Q{mac}=[ 6  0  2 12  0  0  0  0]

        sign=8'b00110000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001001, 8'b00001110, 8'b00011010, 8'b01000010, 8'b00000111, 8'b00011011, 8'b00101111, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00001001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 39: 
        // x=-64, 
        // s=[-1. -1. -1.  1.  1. -1.  1. -1.],
        // w=[16  3 18 15  9  7 12  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  7877.   -832.   4186.  12000.  -1833. -20021.  -6892.  -7405.], 
        // Q{mac}=[ 7  0  4 11  0  0  0  0]

        sign=8'b00011010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00010000, 8'b00000011, 8'b00010010, 8'b00001111, 8'b00001001, 8'b00000111, 8'b00001100, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 40: 
        // x=-91, 
        // s=[-1. -1.  1.  1. -1. -1. -1. -1.],
        // w=[17 23 59  5  9 22  5  4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  9424.   1261.  -1183.  11545.  -1014. -18019.  -6437.  -7041.], 
        // Q{mac}=[ 9  1  0 11  0  0  0  0]

        sign=8'b00110000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00010001, 8'b00010111, 8'b00111011, 8'b00000101, 8'b00001001, 8'b00010110, 8'b00000101, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10100101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 41: 
        // x=118, 
        // s=[-1. -1.  1. -1.  1. -1.  1. -1.],
        // w=[37  2 62 36 10  4  9  7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  5058.   1025.   6133.   7297.    166. -18491.  -5375.  -7867.], 
        // Q{mac}=[4 1 5 7 0 0 0 0]

        sign=8'b00101010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00100101, 8'b00000010, 8'b00111110, 8'b00100100, 8'b00001010, 8'b00000100, 8'b00001001, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b01110110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 42: 
        // x=-37, 
        // s=[ 1.  1. -1. -1.  1. -1. -1.  1.],
        // w=[ 55 125  24   1  34  15 124   2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  3023.  -3600.   7021.   7334.  -1092. -17936.   -787.  -7941.], 
        // Q{mac}=[2 0 6 7 0 0 0 0]

        sign=8'b11001001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00110111, 8'b01111101, 8'b00011000, 8'b00000001, 8'b00100010, 8'b00001111, 8'b01111100, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11011011;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 43: 
        // x=14, 
        // s=[ 1.  1. -1. -1.  1. -1. -1. -1.],
        // w=[10 17  8 11 16  6 16  6],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  3163.  -3362.   6909.   7180.   -868. -18020.  -1011.  -8025.], 
        // Q{mac}=[3 0 6 7 0 0 0 0]

        sign=8'b11001000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001010, 8'b00010001, 8'b00001000, 8'b00001011, 8'b00010000, 8'b00000110, 8'b00010000, 8'b00000110};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00001110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 44: 
        // x=-119, 
        // s=[ 1. -1.  1.  1. -1. -1. -1. -1.],
        // w=[6 4 2 2 9 3 7 5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  2449.  -2886.   6671.   6942.    203. -17663.   -178.  -7430.], 
        // Q{mac}=[2 0 6 6 0 0 0 0]

        sign=8'b10110000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000110, 8'b00000100, 8'b00000010, 8'b00000010, 8'b00001001, 8'b00000011, 8'b00000111, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 45: 
        // x=-120, 
        // s=[-1. -1.  1.  1. -1. -1. -1.  1.],
        // w=[4 8 4 5 1 5 7 9],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  2929.  -1926.   6191.   6342.    323. -17063.    662.  -8510.], 
        // Q{mac}=[2 0 6 6 0 0 0 0]

        sign=8'b00110001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000100, 8'b00001000, 8'b00000100, 8'b00000101, 8'b00000001, 8'b00000101, 8'b00000111, 8'b00001001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 46: 
        // x=-73, 
        // s=[ 1. -1. -1. -1. -1. -1.  1.  1.],
        // w=[11  6  4  2  2  9  3  0],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  2126.  -1488.   6483.   6488.    469. -16406.    443.  -8510.], 
        // Q{mac}=[2 0 6 6 0 0 0 0]

        sign=8'b10000011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001011, 8'b00000110, 8'b00000100, 8'b00000010, 8'b00000010, 8'b00001001, 8'b00000011, 8'b00000000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10110111;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 47: 
        // x=-120, 
        // s=[ 1. -1.  1.  1. -1.  1. -1. -1.],
        // w=[ 6  4  2  8 12  0  7  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  1406.  -1008.   6243.   5528.   1909. -16406.   1283.  -8150.], 
        // Q{mac}=[1 0 6 5 1 0 1 0]

        sign=8'b10110100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000110, 8'b00000100, 8'b00000010, 8'b00001000, 8'b00001100, 8'b00000000, 8'b00000111, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 48: 
        // x=-121, 
        // s=[ 1. -1. -1.  1. -1.  1. -1.  1.],
        // w=[2 8 1 7 1 3 5 4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  1164.    -40.   6364.   4681.   2030. -16769.   1888.  -8634.], 
        // Q{mac}=[1 0 6 4 1 0 1 0]

        sign=8'b10010101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00001000, 8'b00000001, 8'b00000111, 8'b00000001, 8'b00000011, 8'b00000101, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000111;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 49: 
        // x=-78, 
        // s=[-1.  1. -1.  1. -1.  1. -1.  1.],
        // w=[2 1 3 0 2 1 1 8],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  1320.   -118.   6598.   4681.   2186. -16847.   1966.  -9258.], 
        // Q{mac}=[1 0 6 4 2 0 1 0]

        sign=8'b01010101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00000001, 8'b00000011, 8'b00000000, 8'b00000010, 8'b00000001, 8'b00000001, 8'b00001000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10110010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 50: 
        // x=115, 
        // s=[-1. -1.  1. -1.  1.  1.  1. -1.],
        // w=[39  9 69 34  8  1  8  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -3165.  -1153.  14533.    771.   3106. -16732.   2886.  -9603.], 
        // Q{mac}=[ 0  0 14  0  3  0  2  0]

        sign=8'b00101110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00100111, 8'b00001001, 8'b01000101, 8'b00100010, 8'b00001000, 8'b00000001, 8'b00001000, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b01110011;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 51: 
        // x=-37, 
        // s=[ 1.  1. -1.  1.  1. -1. -1. -1.],
        // w=[ 61 118  11   8  32  15 127   6],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -5422.  -5519.  14940.    475.   1922. -16177.   7585.  -9381.], 
        // Q{mac}=[ 0  0 14  0  1  0  7  0]

        sign=8'b11011000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00111101, 8'b01110110, 8'b00001011, 8'b00001000, 8'b00100000, 8'b00001111, 8'b01111111, 8'b00000110};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11011011;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 52: 
        // x=18, 
        // s=[ 1.  1. -1. -1.  1. -1. -1. -1.],
        // w=[ 4 26  9  9  8  7 14  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -5350.  -5051.  14778.    313.   2066. -16303.   7333.  -9435.], 
        // Q{mac}=[ 0  0 14  0  2  0  7  0]

        sign=8'b11001000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000100, 8'b00011010, 8'b00001001, 8'b00001001, 8'b00001000, 8'b00000111, 8'b00001110, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00010010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 53: 
        // x=119, 
        // s=[-1. -1.  1. -1.  1. -1. -1. -1.],
        // w=[41  5 64 34 10  9  1  7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-10229.  -5646.  22394.  -3733.   3256. -17374.   7214. -10268.], 
        // Q{mac}=[ 0  0 21  0  3  0  7  0]

        sign=8'b00101000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00101001, 8'b00000101, 8'b01000000, 8'b00100010, 8'b00001010, 8'b00001001, 8'b00000001, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b01110111;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 54: 
        // x=-34, 
        // s=[ 1.  1. -1.  1.  1. -1. -1. -1.],
        // w=[ 48 114  20   6  36  15 124   1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-11861.  -9522.  23074.  -3937.   2032. -16864.  11430. -10234.], 
        // Q{mac}=[ 0  0 22  0  1  0 11  0]

        sign=8'b11011000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00110000, 8'b01110010, 8'b00010100, 8'b00000110, 8'b00100100, 8'b00001111, 8'b01111100, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11011110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 55: 
        // x=-11, 
        // s=[ 1.  1. -1. -1.  1. -1. -1. -1.],
        // w=[ 4 12  7 17  8  7 17  8],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-11905.  -9654.  23151.  -3750.   1944. -16787.  11617. -10146.], 
        // Q{mac}=[ 0  0 22  0  1  0 11  0]

        sign=8'b11001000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000100, 8'b00001100, 8'b00000111, 8'b00010001, 8'b00001000, 8'b00000111, 8'b00010001, 8'b00001000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11110101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 56: 
        // x=-3, 
        // s=[-1. -1.  1. -1. -1.  1. -1. -1.],
        // w=[23 14 60 31 47 28 15  7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-11836.  -9612.  22971.  -3657.   2085. -16871.  11662. -10125.], 
        // Q{mac}=[ 0  0 22  0  2  0 11  0]

        sign=8'b00100100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00010111, 8'b00001110, 8'b00111100, 8'b00011111, 8'b00101111, 8'b00011100, 8'b00001111, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11111101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 57: 
        // x=105, 
        // s=[-1. -1.  1. -1.  1. -1.  1.  1.],
        // w=[39 15 64 35 16 15 10  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-15931. -11187.  29691.  -7332.   3765. -18446.  12712.  -9810.], 
        // Q{mac}=[ 0  0 28  0  3  0 12  0]

        sign=8'b00101011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00100111, 8'b00001111, 8'b01000000, 8'b00100011, 8'b00010000, 8'b00001111, 8'b00001010, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b01101001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 58: 
        // x=-111, 
        // s=[ 1.  1. -1.  1. -1.  1.  1. -1.],
        // w=[29  4 36 23 19 12  0  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-19150. -11631.  33687.  -9885.   5874. -19778.  12712.  -9255.], 
        // Q{mac}=[ 0  0 32  0  5  0 12  0]

        sign=8'b11010110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00011101, 8'b00000100, 8'b00100100, 8'b00010111, 8'b00010011, 8'b00001100, 8'b00000000, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10010001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 59: 
        // x=-124, 
        // s=[ 1.  1. -1.  1.  1.  1. -1. -1.],
        // w=[29  3 35 23  5  7 18  4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-22746. -12003.  38027. -12737.   5254. -20646.  14944.  -8759.], 
        // Q{mac}=[ 0  0 37  0  5  0 14  0]

        sign=8'b11011100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00011101, 8'b00000011, 8'b00100011, 8'b00010111, 8'b00000101, 8'b00000111, 8'b00010010, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000100;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 60: 
        // x=-122, 
        // s=[-1.  1. -1.  1. -1.  1. -1.  1.],
        // w=[4 4 6 5 5 1 2 6],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-22258. -12491.  38759. -13347.   5864. -20768.  15188.  -9491.], 
        // Q{mac}=[ 0  0 37  0  5  0 14  0]

        sign=8'b01010101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000100, 8'b00000100, 8'b00000110, 8'b00000101, 8'b00000101, 8'b00000001, 8'b00000010, 8'b00000110};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 61: 
        // x=-122, 
        // s=[ 1. -1.  1.  1. -1. -1. -1. -1.],
        // w=[ 2  2  3  0  5 10  1  6],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-22502. -12247.  38393. -13347.   6474. -19548.  15310.  -8759.], 
        // Q{mac}=[ 0  0 37  0  6  0 14  0]

        sign=8'b10110000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00000010, 8'b00000011, 8'b00000000, 8'b00000101, 8'b00001010, 8'b00000001, 8'b00000110};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 62: 
        // x=-98, 
        // s=[ 1.  1. -1.  1. -1.  1.  1.  1.],
        // w=[ 4  1  8  0 13  3  1  0],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-22894. -12345.  39177. -13347.   7748. -19842.  15212.  -8759.], 
        // Q{mac}=[ 0  0 38  0  7  0 14  0]

        sign=8'b11010111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000100, 8'b00000001, 8'b00001000, 8'b00000000, 8'b00001101, 8'b00000011, 8'b00000001, 8'b00000000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10011110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 63: 
        // x=-55, 
        // s=[ 1.  1. -1. -1. -1.  1.  1.  1.],
        // w=[11  7 18 15 34 40  4  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-23499. -12730.  40167. -12522.   9618. -22042.  14992.  -8924.], 
        // Q{mac}=[ 0  0 39  0  9  0 14  0]

        sign=8'b11000111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001011, 8'b00000111, 8'b00010010, 8'b00001111, 8'b00100010, 8'b00101000, 8'b00000100, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11001001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 64: 
        // x=-128, 
        // s=[ 1.  1.  1.  1. -1.  1. -1. -1.],
        // w=[18 18 14  1  8 15 24  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-25803. -15034.  38375. -12650.  10642. -23962.  18064.  -8284.], 
        // Q{mac}=[ 0  0 37  0 10  0 17  0]

        sign=8'b11110100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00010010, 8'b00010010, 8'b00001110, 8'b00000001, 8'b00001000, 8'b00001111, 8'b00011000, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 65: 
        // x=27, 
        // s=[-1. -1. -1.  1.  1. -1.  1. -1.],
        // w=[18 13  2 11  7 16  3  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-26289. -15385.  38321. -12353.  10831. -24394.  18145.  -8419.], 
        // Q{mac}=[ 0  0 37  0 10  0 17  0]

        sign=8'b00011010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00010010, 8'b00001101, 8'b00000010, 8'b00001011, 8'b00000111, 8'b00010000, 8'b00000011, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00011011;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 66: 
        // x=-56, 
        // s=[-1. -1.  1.  1.  1. -1. -1.  1.],
        // w=[ 2  9 18 14  0 16 12  7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-26177. -14881.  37313. -13137.  10831. -23498.  18817.  -8811.], 
        // Q{mac}=[ 0  0 36  0 10  0 18  0]

        sign=8'b00111001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00001001, 8'b00010010, 8'b00001110, 8'b00000000, 8'b00010000, 8'b00001100, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11001000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 67: 
        // x=54, 
        // s=[ 1.  1. -1. -1.  1.  1.  1.  1.],
        // w=[ 8 15  6 15  5  2  5  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-25745. -14071.  36989. -13947.  11101. -23390.  19087.  -8649.], 
        // Q{mac}=[ 0  0 36  0 10  0 18  0]

        sign=8'b11001111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001000, 8'b00001111, 8'b00000110, 8'b00001111, 8'b00000101, 8'b00000010, 8'b00000101, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00110110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 68: 
        // x=-56, 
        // s=[-1. -1.  1.  1. -1. -1. -1.  1.],
        // w=[ 4  7  9  9 13 10 12  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-25521. -13679.  36485. -14451.  11829. -22830.  19759.  -8761.], 
        // Q{mac}=[ 0  0 35  0 11  0 19  0]

        sign=8'b00110001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000100, 8'b00000111, 8'b00001001, 8'b00001001, 8'b00001101, 8'b00001010, 8'b00001100, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11001000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 69: 
        // x=54, 
        // s=[-1.  1. -1.  1.  1.  1.  1. -1.],
        // w=[ 6  8  5  0 13  8 12  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-25845. -13247.  36215. -14451.  12531. -22398.  20407.  -8869.], 
        // Q{mac}=[ 0  0 35  0 12  0 19  0]

        sign=8'b01011110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000110, 8'b00001000, 8'b00000101, 8'b00000000, 8'b00001101, 8'b00001000, 8'b00001100, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00110110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 70: 
        // x=-102, 
        // s=[-1. -1. -1. -1.  1. -1. -1. -1.],
        // w=[12  4  5  2 29 21  9  4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-24621. -12839.  36725. -14247.   9573. -20256.  21325.  -8461.], 
        // Q{mac}=[ 0  0 35  0  9  0 20  0]

        sign=8'b00001000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001100, 8'b00000100, 8'b00000101, 8'b00000010, 8'b00011101, 8'b00010101, 8'b00001001, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10011010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 71: 
        // x=99, 
        // s=[ 1. -1.  1. -1. -1.  1.  1. -1.],
        // w=[ 2  6  0  6 25 26 13 10],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-24423. -13433.  36725. -14841.   7098. -17682.  22612.  -9451.], 
        // Q{mac}=[ 0  0 35  0  6  0 22  0]

        sign=8'b10100110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00000110, 8'b00000000, 8'b00000110, 8'b00011001, 8'b00011010, 8'b00001101, 8'b00001010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b01100011;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 72: 
        // x=-100, 
        // s=[-1. -1. -1.  1.  1. -1. -1.  1.],
        // w=[12  2  1  8 21 24 13  4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-23223. -13233.  36825. -15641.   4998. -15282.  23912.  -9851.], 
        // Q{mac}=[ 0  0 35  0  4  0 23  0]

        sign=8'b00011001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001100, 8'b00000010, 8'b00000001, 8'b00001000, 8'b00010101, 8'b00011000, 8'b00001101, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10011100;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 73: 
        // x=99, 
        // s=[ 1. -1.  1. -1. -1.  1.  1. -1.],
        // w=[ 6  1  8  7 20 18  5  6],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-22629. -13332.  37617. -16334.   3018. -13500.  24407. -10445.], 
        // Q{mac}=[ 0  0 36  0  2  0 23  0]

        sign=8'b10100110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000110, 8'b00000001, 8'b00001000, 8'b00000111, 8'b00010100, 8'b00010010, 8'b00000101, 8'b00000110};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b01100011;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 74: 
        // x=-127, 
        // s=[-1.  1. -1.  1.  1. -1. -1.  1.],
        // w=[ 2  1  7  5  8 20 10  4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-22375. -13459.  38506. -16969.   2002. -10960.  25677. -10953.], 
        // Q{mac}=[ 0  0 37  0  1  0 25  0]

        sign=8'b01011001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00000001, 8'b00000111, 8'b00000101, 8'b00001000, 8'b00010100, 8'b00001010, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 75: 
        // x=125, 
        // s=[ 1.  1.  1. -1. -1.  1.  1. -1.],
        // w=[ 3  0 14  4 15  5  3 12],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-22000. -13459.  40256. -17469.    127. -10335.  26052. -12453.], 
        // Q{mac}=[ 0  0 39  0  0  0 25  0]

        sign=8'b11100110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00000000, 8'b00001110, 8'b00000100, 8'b00001111, 8'b00000101, 8'b00000011, 8'b00001100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b01111101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 76: 
        // x=-127, 
        // s=[-1. -1. -1.  1.  1. -1.  1. -1.],
        // w=[10  1 18  2 12 17  2  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-20730. -13332.  42542. -17723.  -1397.  -8176.  25798. -12199.], 
        // Q{mac}=[ 0  0 41  0  0  0 25  0]

        sign=8'b00011010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001010, 8'b00000001, 8'b00010010, 8'b00000010, 8'b00001100, 8'b00010001, 8'b00000010, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 77: 
        // x=125, 
        // s=[ 1. -1.  1. -1. -1.  1. -1. -1.],
        // w=[ 7  4 10  1  3 13  3  7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-19855. -13832.  43792. -17848.  -1772.  -6551.  25423. -13074.], 
        // Q{mac}=[ 0  0 42  0  0  0 24  0]

        sign=8'b10100100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00000100, 8'b00001010, 8'b00000001, 8'b00000011, 8'b00001101, 8'b00000011, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b01111101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 78: 
        // x=124, 
        // s=[ 1.  1. -1.  1. -1.  1.  1.  1.],
        // w=[ 9 11 11 11  4  5  9  0],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-18739. -12468.  42428. -16484.  -2268.  -5931.  26539. -13074.], 
        // Q{mac}=[ 0  0 41  0  0  0 25  0]

        sign=8'b11010111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001001, 8'b00001011, 8'b00001011, 8'b00001011, 8'b00000100, 8'b00000101, 8'b00001001, 8'b00000000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b01111100;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 79: 
        // x=-128, 
        // s=[ 1. -1.  1.  1. -1.  1. -1. -1.],
        // w=[ 6  7  9 21  9 15  7  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-19507. -11572.  41276. -19172.  -1116.  -7851.  27435. -12434.], 
        // Q{mac}=[ 0  0 40  0  0  0 26  0]

        sign=8'b10110100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000110, 8'b00000111, 8'b00001001, 8'b00010101, 8'b00001001, 8'b00001111, 8'b00000111, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 80: 
        // x=-123, 
        // s=[-1.  1.  1. -1. -1. -1.  1. -1.],
        // w=[ 1  5  7 16  4  7  0  8],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-19384. -12187.  40415. -17204.   -624.  -6990.  27435. -11450.], 
        // Q{mac}=[ 0  0 39  0  0  0 26  0]

        sign=8'b01100010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00000101, 8'b00000111, 8'b00010000, 8'b00000100, 8'b00000111, 8'b00000000, 8'b00001000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 81: 
        // x=8, 
        // s=[-1. -1.  1.  1.  1. -1.  1. -1.],
        // w=[ 7  2  2  9 13 10  2  9],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-19440. -12203.  40431. -17132.   -520.  -7070.  27451. -11522.], 
        // Q{mac}=[ 0  0 39  0  0  0 26  0]

        sign=8'b00111010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00000010, 8'b00000010, 8'b00001001, 8'b00001101, 8'b00001010, 8'b00000010, 8'b00001001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00001000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 82: 
        // x=5, 
        // s=[-1.  1. -1.  1. -1.  1.  1.  1.],
        // w=[ 6  2  6  0  8 16  6  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-19470. -12193.  40401. -17132.   -560.  -6990.  27481. -11507.], 
        // Q{mac}=[ 0  0 39  0  0  0 26  0]

        sign=8'b01010111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000110, 8'b00000010, 8'b00000110, 8'b00000000, 8'b00001000, 8'b00010000, 8'b00000110, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00000101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 83: 
        // x=-15, 
        // s=[-1.  1.  1.  1. -1. -1. -1.  1.],
        // w=[ 3  5  8 14  2  5  5 10],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-19425. -12268.  40281. -17342.   -530.  -6915.  27556. -11657.], 
        // Q{mac}=[ 0  0 39  0  0  0 26  0]

        sign=8'b01110001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00000101, 8'b00001000, 8'b00001110, 8'b00000010, 8'b00000101, 8'b00000101, 8'b00001010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11110001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 84: 
        // x=-117, 
        // s=[-1.  1. -1. -1.  1.  1.  1. -1.],
        // w=[5 9 2 4 1 5 3 2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-18840. -13321.  40515. -16874.   -647.  -7500.  27205. -11423.], 
        // Q{mac}=[ 0  0 39  0  0  0 26  0]

        sign=8'b01001110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000101, 8'b00001001, 8'b00000010, 8'b00000100, 8'b00000001, 8'b00000101, 8'b00000011, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001011;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 85: 
        // x=-121, 
        // s=[-1. -1.  1. -1.  1. -1. -1.  1.],
        // w=[ 3  6 11  6  9  4  5  7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-18477. -12595.  39184. -16148.  -1736.  -7016.  27810. -12270.], 
        // Q{mac}=[ 0  0 38  0  0  0 27  0]

        sign=8'b00101001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00000110, 8'b00001011, 8'b00000110, 8'b00001001, 8'b00000100, 8'b00000101, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000111;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 86: 
        // x=-120, 
        // s=[ 1.  1.  1. -1.  1. -1. -1. -1.],
        // w=[ 0  3  2  9 14  5  4  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-18477. -12955.  38944. -15068.  -3416.  -6416.  28290. -12030.], 
        // Q{mac}=[ 0  0 38  0  0  0 27  0]

        sign=8'b11101000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000000, 8'b00000011, 8'b00000010, 8'b00001001, 8'b00001110, 8'b00000101, 8'b00000100, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 87: 
        // x=-118, 
        // s=[-1.  1. -1. -1.  1.  1.  1.  1.],
        // w=[3 3 3 5 8 8 7 1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-18123. -13309.  39298. -14478.  -4360.  -7360.  27464. -12148.], 
        // Q{mac}=[ 0  0 38  0  0  0 26  0]

        sign=8'b01001111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00000011, 8'b00000011, 8'b00000101, 8'b00001000, 8'b00001000, 8'b00000111, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 88: 
        // x=-120, 
        // s=[-1. -1.  1. -1.  1. -1.  1.  1.],
        // w=[14  3  1  2 11  6  0 10],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-16443. -12949.  39178. -14238.  -5680.  -6640.  27464. -13348.], 
        // Q{mac}=[ 0  0 38  0  0  0 26  0]

        sign=8'b00101011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001110, 8'b00000011, 8'b00000001, 8'b00000010, 8'b00001011, 8'b00000110, 8'b00000000, 8'b00001010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 89: 
        // x=-122, 
        // s=[-1. -1.  1. -1.  1. -1. -1. -1.],
        // w=[ 1  5  4  7 12  7 10  4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-16321. -12339.  38690. -13384.  -7144.  -5786.  28684. -12860.], 
        // Q{mac}=[ 0  0 37  0  0  0 28  0]

        sign=8'b00101000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00000101, 8'b00000100, 8'b00000111, 8'b00001100, 8'b00000111, 8'b00001010, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 90: 
        // x=-116, 
        // s=[ 1.  1. -1. -1.  1. -1.  1.  1.],
        // w=[ 7 15 20 14 20  1  1  0],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-17133. -14079.  41010. -11760.  -9464.  -5670.  28568. -12860.], 
        // Q{mac}=[ 0  0 40  0  0  0 27  0]

        sign=8'b11001011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00001111, 8'b00010100, 8'b00001110, 8'b00010100, 8'b00000001, 8'b00000001, 8'b00000000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001100;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 91: 
        // x=-122, 
        // s=[-1.  1. -1.  1.  1. -1. -1.  1.],
        // w=[ 3 12  6  0 12  9  6 10],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-16767. -15543.  41742. -11760. -10928.  -4572.  29300. -14080.], 
        // Q{mac}=[ 0  0 40  0  0  0 28  0]

        sign=8'b01011001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00001100, 8'b00000110, 8'b00000000, 8'b00001100, 8'b00001001, 8'b00000110, 8'b00001010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 92: 
        // x=-115, 
        // s=[ 1.  1. -1. -1.  1. -1.  1. -1.],
        // w=[ 3  4 12 12 10  9  2  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-17112. -16003.  43122. -10380. -12078.  -3537.  29070. -13735.], 
        // Q{mac}=[ 0  0 42  0  0  0 28  0]

        sign=8'b11001010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00000100, 8'b00001100, 8'b00001100, 8'b00001010, 8'b00001001, 8'b00000010, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 93: 
        // x=114, 
        // s=[ 1.  1. -1.  1.  1. -1. -1. -1.],
        // w=[12 18 10  5 29 27  1  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-15744. -13951.  41982.  -9810.  -8772.  -6615.  28956. -13963.], 
        // Q{mac}=[ 0  0 40  0  0  0 28  0]

        sign=8'b11011000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001100, 8'b00010010, 8'b00001010, 8'b00000101, 8'b00011101, 8'b00011011, 8'b00000001, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b01110010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 94: 
        // x=120, 
        // s=[ 1.  1. -1.  1.  1. -1.  1. -1.],
        // w=[11  3 12  1  5  1  6  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-14424. -13591.  40542.  -9690.  -8172.  -6735.  29676. -14563.], 
        // Q{mac}=[ 0  0 39  0  0  0 28  0]

        sign=8'b11011010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001011, 8'b00000011, 8'b00001100, 8'b00000001, 8'b00000101, 8'b00000001, 8'b00000110, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b01111000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 95: 
        // x=120, 
        // s=[ 1.  1. -1.  1. -1.  1.  1. -1.],
        // w=[15  4  6  5 19 13  3  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-12624. -13111.  39822.  -9090. -10452.  -5175.  30036. -14803.], 
        // Q{mac}=[ 0  0 38  0  0  0 29  0]

        sign=8'b11010110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001111, 8'b00000100, 8'b00000110, 8'b00000101, 8'b00010011, 8'b00001101, 8'b00000011, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b01111000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 96: 
        // x=-120, 
        // s=[-1. -1. -1.  1.  1. -1. -1. -1.],
        // w=[ 9  8  4  2 13  4  4  4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-11544. -12151.  40302.  -9330. -12012.  -4695.  30516. -14323.], 
        // Q{mac}=[ 0  0 39  0  0  0 29  0]

        sign=8'b00011000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001001, 8'b00001000, 8'b00000100, 8'b00000010, 8'b00001101, 8'b00000100, 8'b00000100, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 97: 
        // x=-128, 
        // s=[-1.  1.  1.  1.  1.  1. -1. -1.],
        // w=[7 2 2 0 2 2 4 2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-10648. -12407.  40046.  -9330. -12268.  -4951.  31028. -14067.], 
        // Q{mac}=[ 0  0 39  0  0  0 30  0]

        sign=8'b01111100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00000010, 8'b00000010, 8'b00000000, 8'b00000010, 8'b00000010, 8'b00000100, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 98: 
        // x=-128, 
        // s=[-1.  1.  1. -1.  1.  1.  1.  1.],
        // w=[7 0 4 4 5 0 2 9],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -9752. -12407.  39534.  -8818. -12908.  -4951.  30772. -15219.], 
        // Q{mac}=[ 0  0 38  0  0  0 30  0]

        sign=8'b01101111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00000000, 8'b00000100, 8'b00000100, 8'b00000101, 8'b00000000, 8'b00000010, 8'b00001001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 99: 
        // x=-128, 
        // s=[ 1. -1. -1. -1.  1. -1.  1.  1.],
        // w=[3 5 5 7 4 8 5 7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-10136. -11767.  40174.  -7922. -13420.  -3927.  30132. -16115.], 
        // Q{mac}=[ 0  0 39  0  0  0 29  0]

        sign=8'b10001011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00000101, 8'b00000101, 8'b00000111, 8'b00000100, 8'b00001000, 8'b00000101, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 100: 
        // x=-120, 
        // s=[ 1. -1.  1. -1. -1.  1.  1.  1.],
        // w=[2 2 5 8 3 4 6 4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[-10376. -11527.  39574.  -6962. -13060.  -4407.  29412. -16595.], 
        // Q{mac}=[ 0  0 38  0  0  0 28  0]

        sign=8'b10100111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00000010, 8'b00000101, 8'b00001000, 8'b00000011, 8'b00000100, 8'b00000110, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 101: 
        // x=-122, 
        // s=[-1. -1.  1. -1.  1.  1.  1.  1.],
        // w=[ 7 13  8  3  3  3  3  1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -9522.  -9941.  38598.  -6596. -13426.  -4773.  29046. -16717.], 
        // Q{mac}=[ 0  0 37  0  0  0 28  0]

        sign=8'b00101111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00001101, 8'b00001000, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 102: 
        // x=-125, 
        // s=[-1. -1.  1.  1.  1.  1. -1. -1.],
        // w=[ 8  7  5  0 13  1  8  4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -8522.  -9066.  37973.  -6596. -15051.  -4898.  30046. -16217.], 
        // Q{mac}=[ 0  0 37  0  0  0 29  0]

        sign=8'b00111100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001000, 8'b00000111, 8'b00000101, 8'b00000000, 8'b00001101, 8'b00000001, 8'b00001000, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000011;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 103: 
        // x=-12, 
        // s=[-1. -1.  1.  1.  1.  1.  1. -1.],
        // w=[ 6  2 11  2 12 12  6  4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -8450.  -9042.  37841.  -6620. -15195.  -5042.  29974. -16169.], 
        // Q{mac}=[ 0  0 36  0  0  0 29  0]

        sign=8'b00111110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000110, 8'b00000010, 8'b00001011, 8'b00000010, 8'b00001100, 8'b00001100, 8'b00000110, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11110100;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 104: 
        // x=-41, 
        // s=[-1. -1.  1. -1.  1.  1.  1. -1.],
        // w=[ 8  4  9  1 12  5 11  8],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -8122.  -8878.  37472.  -6579. -15687.  -5247.  29523. -15841.], 
        // Q{mac}=[ 0  0 36  0  0  0 28  0]

        sign=8'b00101110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001000, 8'b00000100, 8'b00001001, 8'b00000001, 8'b00001100, 8'b00000101, 8'b00001011, 8'b00001000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11010111;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 105: 
        // x=-66, 
        // s=[-1. -1.  1. -1.  1.  1. -1. -1.],
        // w=[ 5  3 19  1 18  7 12  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -7792.  -8680.  36218.  -6513. -16875.  -5709.  30315. -15709.], 
        // Q{mac}=[ 0  0 35  0  0  0 29  0]

        sign=8'b00101100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000101, 8'b00000011, 8'b00010011, 8'b00000001, 8'b00010010, 8'b00000111, 8'b00001100, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10111110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 106: 
        // x=65, 
        // s=[-1. -1. -1.  1. -1. -1.  1.  1.],
        // w=[ 2  6 10  7 10  4 15  1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -7922.  -9070.  35568.  -6058. -17525.  -5969.  31290. -15644.], 
        // Q{mac}=[ 0  0 34  0  0  0 30  0]

        sign=8'b00010011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00000110, 8'b00001010, 8'b00000111, 8'b00001010, 8'b00000100, 8'b00001111, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b01000001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 107: 
        // x=-30, 
        // s=[-1. -1.  1.  1. -1. -1.  1.  1.],
        // w=[18 25 38 19 16  4  3  6],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -7382.  -8320.  34428.  -6628. -17045.  -5849.  31200. -15824.], 
        // Q{mac}=[ 0  0 33  0  0  0 30  0]

        sign=8'b00110011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00010010, 8'b00011001, 8'b00100110, 8'b00010011, 8'b00010000, 8'b00000100, 8'b00000011, 8'b00000110};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11100010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 108: 
        // x=62, 
        // s=[-1. -1.  1.  1.  1. -1. -1. -1.],
        // w=[10  9  5 19  0  6  2  7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -8002.  -8878.  34738.  -5450. -17045.  -6221.  31076. -16258.], 
        // Q{mac}=[ 0  0 33  0  0  0 30  0]

        sign=8'b00111000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001010, 8'b00001001, 8'b00000101, 8'b00010011, 8'b00000000, 8'b00000110, 8'b00000010, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00111110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 109: 
        // x=39, 
        // s=[-1. -1.  1.  1.  1. -1. -1.  1.],
        // w=[15 12 34 32  2 11  6  4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -8587.  -9346.  36064.  -4202. -16967.  -6650.  30842. -16102.], 
        // Q{mac}=[ 0  0 35  0  0  0 30  0]

        sign=8'b00111001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001111, 8'b00001100, 8'b00100010, 8'b00100000, 8'b00000010, 8'b00001011, 8'b00000110, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00100111;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 110: 
        // x=28, 
        // s=[-1. -1. -1.  1. -1. -1.  1. -1.],
        // w=[ 3  6 20  1  4  7 26  1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -8671.  -9514.  35504.  -4174. -17079.  -6846.  31570. -16130.], 
        // Q{mac}=[ 0  0 34  0  0  0 30  0]

        sign=8'b00010010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00000110, 8'b00010100, 8'b00000001, 8'b00000100, 8'b00000111, 8'b00011010, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00011100;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 111: 
        // x=14, 
        // s=[-1. -1. -1.  1. -1. -1.  1.  1.],
        // w=[13  7 14 17  4  6 23  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -8853.  -9612.  35308.  -3936. -17135.  -6930.  31892. -16060.], 
        // Q{mac}=[ 0  0 34  0  0  0 31  0]

        sign=8'b00010011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001101, 8'b00000111, 8'b00001110, 8'b00010001, 8'b00000100, 8'b00000110, 8'b00010111, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00001110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 112: 
        // x=27, 
        // s=[ 1.  1.  1.  1. -1.  1. -1. -1.],
        // w=[ 5  6  4  0  5  5 13 13],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -8718.  -9450.  35416.  -3936. -17270.  -6795.  31541. -16411.], 
        // Q{mac}=[ 0  0 34  0  0  0 30  0]

        sign=8'b11110100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000101, 8'b00000110, 8'b00000100, 8'b00000000, 8'b00000101, 8'b00000101, 8'b00001101, 8'b00001101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00011011;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 113: 
        // x=53, 
        // s=[-1. -1. -1.  1.  1. -1.  1. -1.],
        // w=[16 17  7 11 12 13 18  6],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -9566. -10351.  35045.  -3353. -16634.  -7484.  32495. -16729.], 
        // Q{mac}=[ 0  0 34  0  0  0 31  0]

        sign=8'b00011010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00010000, 8'b00010001, 8'b00000111, 8'b00001011, 8'b00001100, 8'b00001101, 8'b00010010, 8'b00000110};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00110101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 114: 
        // x=-12, 
        // s=[ 1. -1.  1.  1.  1. -1.  1. -1.],
        // w=[ 1 13  1 11  7 19 16  4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -9578. -10195.  35033.  -3485. -16718.  -7256.  32303. -16681.], 
        // Q{mac}=[ 0  0 34  0  0  0 31  0]

        sign=8'b10111010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00001101, 8'b00000001, 8'b00001011, 8'b00000111, 8'b00010011, 8'b00010000, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11110100;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 115: 
        // x=17, 
        // s=[-1. -1. -1.  1.  1. -1.  1.  1.],
        // w=[16 17 24 14 30 37 22 11],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -9850. -10484.  34625.  -3247. -16208.  -7885.  32677. -16494.], 
        // Q{mac}=[ 0  0 33  0  0  0 31  0]

        sign=8'b00011011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00010000, 8'b00010001, 8'b00011000, 8'b00001110, 8'b00011110, 8'b00100101, 8'b00010110, 8'b00001011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00010001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 116: 
        // x=-26, 
        // s=[-1. -1. -1.  1.  1. -1.  1.  1.],
        // w=[20 13 28  7 22 23 23  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -9330. -10146.  35353.  -3429. -16780.  -7287.  32079. -16624.], 
        // Q{mac}=[ 0  0 34  0  0  0 31  0]

        sign=8'b00011011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00010100, 8'b00001101, 8'b00011100, 8'b00000111, 8'b00010110, 8'b00010111, 8'b00010111, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11100110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 117: 
        // x=8, 
        // s=[-1.  1. -1.  1.  1.  1.  1.  1.],
        // w=[17 12  9 10  3 16  7  0],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -9466. -10050.  35281.  -3349. -16756.  -7159.  32135. -16624.], 
        // Q{mac}=[ 0  0 34  0  0  0 31  0]

        sign=8'b01011111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00010001, 8'b00001100, 8'b00001001, 8'b00001010, 8'b00000011, 8'b00010000, 8'b00000111, 8'b00000000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00001000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 118: 
        // x=-35, 
        // s=[-1. -1.  1.  1.  1. -1. -1. -1.],
        // w=[42 12 22 43 31 28 45  9],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -7996.  -9630.  34511.  -4854. -17841.  -6179.  33710. -16309.], 
        // Q{mac}=[ 0  0 33  0  0  0 32  0]

        sign=8'b00111000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00101010, 8'b00001100, 8'b00010110, 8'b00101011, 8'b00011111, 8'b00011100, 8'b00101101, 8'b00001001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11011101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 119: 
        // x=4, 
        // s=[-1.  1.  1.  1.  1. -1. -1. -1.],
        // w=[10 21  0 16 64 21 51  7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -8036.  -9546.  34511.  -4790. -17585.  -6263.  33506. -16337.], 
        // Q{mac}=[ 0  0 33  0  0  0 32  0]

        sign=8'b01111000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001010, 8'b00010101, 8'b00000000, 8'b00010000, 8'b01000000, 8'b00010101, 8'b00110011, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00000100;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 120: 
        // x=-46, 
        // s=[ 1. -1.  1.  1. -1. -1. -1.  1.],
        // w=[24 10 27 26 14  6 25  9],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -9140.  -9086.  33269.  -5986. -16941.  -5987.  34656. -16751.], 
        // Q{mac}=[ 0  0 32  0  0  0 33  0]

        sign=8'b10110001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00011000, 8'b00001010, 8'b00011011, 8'b00011010, 8'b00001110, 8'b00000110, 8'b00011001, 8'b00001001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11010010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 121: 
        // x=14, 
        // s=[ 1. -1. -1. -1.  1. -1.  1.  1.],
        // w=[ 6 12 14  7  3  8 17  6],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -9056.  -9254.  33073.  -6084. -16899.  -6099.  34894. -16667.], 
        // Q{mac}=[ 0  0 32  0  0  0 34  0]

        sign=8'b10001011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000110, 8'b00001100, 8'b00001110, 8'b00000111, 8'b00000011, 8'b00001000, 8'b00010001, 8'b00000110};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00001110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 122: 
        // x=-13, 
        // s=[-1. -1.  1.  1. -1. -1.  1.  1.],
        // w=[23 18 14 16  4 23 14  8],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -8757.  -9020.  32891.  -6292. -16847.  -5800.  34712. -16771.], 
        // Q{mac}=[ 0  0 32  0  0  0 33  0]

        sign=8'b00110011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00010111, 8'b00010010, 8'b00001110, 8'b00010000, 8'b00000100, 8'b00010111, 8'b00001110, 8'b00001000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11110011;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 123: 
        // x=23, 
        // s=[-1.  1. -1. -1. -1.  1.  1. -1.],
        // w=[ 1  4 16 15  5 17 24  6],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -8780.  -8928.  32523.  -6637. -16962.  -5409.  35264. -16909.], 
        // Q{mac}=[ 0  0 31  0  0  0 34  0]

        sign=8'b01000110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00000100, 8'b00010000, 8'b00001111, 8'b00000101, 8'b00010001, 8'b00011000, 8'b00000110};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00010111;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 124: 
        // x=-114, 
        // s=[ 1.  1.  1. -1.  1. -1.  1.  1.],
        // w=[ 3  1  1  6  7  7 10  8],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -9122.  -9042.  32409.  -5953. -17760.  -4611.  34124. -17821.], 
        // Q{mac}=[ 0  0 31  0  0  0 33  0]

        sign=8'b11101011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00000001, 8'b00000001, 8'b00000110, 8'b00000111, 8'b00000111, 8'b00001010, 8'b00001000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 125: 
        // x=-105, 
        // s=[-1. -1.  1.  1.  1.  1. -1.  1.],
        // w=[8 2 3 2 8 5 5 2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -8282.  -8832.  32094.  -6163. -18600.  -5136.  34649. -18031.], 
        // Q{mac}=[ 0  0 31  0  0  0 33  0]

        sign=8'b00111101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001000, 8'b00000010, 8'b00000011, 8'b00000010, 8'b00001000, 8'b00000101, 8'b00000101, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10010111;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 126: 
        // x=-121, 
        // s=[-1. -1.  1.  1. -1.  1. -1.  1.],
        // w=[13  5 10  2  5  3  5  7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -6709.  -8227.  30884.  -6405. -17995.  -5499.  35254. -18878.], 
        // Q{mac}=[ 0  0 30  0  0  0 34  0]

        sign=8'b00110101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001101, 8'b00000101, 8'b00001010, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000101, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000111;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 127: 
        // x=-114, 
        // s=[ 1. -1.  1. -1.  1. -1. -1.  1.],
        // w=[ 2  9  2 14  2 11  3  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -6937.  -7201.  30656.  -4809. -18223.  -4245.  35596. -19106.], 
        // Q{mac}=[ 0  0 29  0  0  0 34  0]

        sign=8'b10101001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00001001, 8'b00000010, 8'b00001110, 8'b00000010, 8'b00001011, 8'b00000011, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 128: 
        // x=-110, 
        // s=[-1. -1.  1. -1. -1.  1. -1.  1.],
        // w=[10  6  5  4  2  3  4  9],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -5837.  -6541.  30106.  -4369. -18003.  -4575.  36036. -20096.], 
        // Q{mac}=[ 0  0 29  0  0  0 35  0]

        sign=8'b00100101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001010, 8'b00000110, 8'b00000101, 8'b00000100, 8'b00000010, 8'b00000011, 8'b00000100, 8'b00001001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10010010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 129: 
        // x=-122, 
        // s=[ 1. -1. -1. -1. -1.  1. -1.  1.],
        // w=[ 1  6  1 12 11 21  3  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -5959.  -5809.  30228.  -2905. -16661.  -7137.  36402. -20462.], 
        // Q{mac}=[ 0  0 29  0  0  0 35  0]

        sign=8'b10000101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00000110, 8'b00000001, 8'b00001100, 8'b00001011, 8'b00010101, 8'b00000011, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 130: 
        // x=-86, 
        // s=[-1. -1.  1. -1. -1.  1.  1. -1.],
        // w=[ 1  6  2 10  3  4  3  1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -5873.  -5293.  30056.  -2045. -16403.  -7481.  36144. -20376.], 
        // Q{mac}=[ 0  0 29  0  0  0 35  0]

        sign=8'b00100110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00000110, 8'b00000010, 8'b00001010, 8'b00000011, 8'b00000100, 8'b00000011, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10101010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 131: 
        // x=-92, 
        // s=[-1.  1.  1. -1.  1. -1. -1.  1.],
        // w=[ 4  1  5  1  2  3 10  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -5505.  -5385.  29596.  -1953. -16587.  -7205.  37064. -20836.], 
        // Q{mac}=[ 0  0 28  0  0  0 36  0]

        sign=8'b01101001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000100, 8'b00000001, 8'b00000101, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00001010, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10100100;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 132: 
        // x=-84, 
        // s=[-1. -1.  1.  1. -1.  1.  1. -1.],
        // w=[ 8  8  6  1  7 12  4  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -4833.  -4713.  29092.  -2037. -15999.  -8213.  36728. -20668.], 
        // Q{mac}=[ 0  0 28  0  0  0 35  0]

        sign=8'b00110110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001000, 8'b00001000, 8'b00000110, 8'b00000001, 8'b00000111, 8'b00001100, 8'b00000100, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10101100;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 133: 
        // x=106, 
        // s=[ 1. -1.  1.  1.  1. -1. -1. -1.],
        // w=[ 4  6 13  9  0  1  5  9],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -4409.  -5349.  30470.  -1083. -15999.  -8319.  36198. -21622.], 
        // Q{mac}=[ 0  0 29  0  0  0 35  0]

        sign=8'b10111000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000100, 8'b00000110, 8'b00001101, 8'b00001001, 8'b00000000, 8'b00000001, 8'b00000101, 8'b00001001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b01101010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 134: 
        // x=104, 
        // s=[ 1.  1. -1.  1. -1. -1.  1.  1.],
        // w=[ 7  7  3  1  3 10  4  0],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -3681.  -4621.  30158.   -979. -16311.  -9359.  36614. -21622.], 
        // Q{mac}=[ 0  0 29  0  0  0 35  0]

        sign=8'b11010011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00000111, 8'b00000011, 8'b00000001, 8'b00000011, 8'b00001010, 8'b00000100, 8'b00000000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b01101000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 135: 
        // x=102, 
        // s=[ 1. -1. -1.  1. -1.  1.  1.  1.],
        // w=[10  3  1  5 24  8  0  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -2661.  -4927.  30056.   -469. -18759.  -8543.  36614. -21316.], 
        // Q{mac}=[ 0  0 29  0  0  0 35  0]

        sign=8'b10010111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001010, 8'b00000011, 8'b00000001, 8'b00000101, 8'b00011000, 8'b00001000, 8'b00000000, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b01100110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 136: 
        // x=-103, 
        // s=[-1. -1. -1. -1.  1.  1.  1. -1.],
        // w=[4 5 6 4 7 4 2 2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -2249.  -4412.  30674.    -57. -19480.  -8955.  36408. -21110.], 
        // Q{mac}=[ 0  0 29  0  0  0 35  0]

        sign=8'b00001110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000100, 8'b00000101, 8'b00000110, 8'b00000100, 8'b00000111, 8'b00000100, 8'b00000010, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10011001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 137: 
        // x=-126, 
        // s=[-1.  1. -1. -1.  1.  1.  1.  1.],
        // w=[1 1 4 6 1 7 1 0],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -2123.  -4538.  31178.    699. -19606.  -9837.  36282. -21110.], 
        // Q{mac}=[ 0  0 30  0  0  0 35  0]

        sign=8'b01001111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00000001, 8'b00000100, 8'b00000110, 8'b00000001, 8'b00000111, 8'b00000001, 8'b00000000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 138: 
        // x=-126, 
        // s=[-1. -1. -1. -1. -1. -1. -1. -1.],
        // w=[3 2 2 2 8 8 8 1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -1745.  -4286.  31430.    951. -18598.  -8829.  37290. -20984.], 
        // Q{mac}=[ 0  0 30  0  0  0 36  0]

        sign=8'b00000000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00001000, 8'b00001000, 8'b00001000, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 139: 
        // x=-128, 
        // s=[ 1. -1. -1. -1. -1. -1. -1.  1.],
        // w=[6 5 5 7 2 1 1 2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -2513.  -3646.  32070.   1847. -18342.  -8701.  37418. -21240.], 
        // Q{mac}=[ 0  0 31  1  0  0 36  0]

        sign=8'b10000001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000110, 8'b00000101, 8'b00000101, 8'b00000111, 8'b00000010, 8'b00000001, 8'b00000001, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 140: 
        // x=-114, 
        // s=[ 1. -1. -1.  1.  1. -1. -1.  1.],
        // w=[ 2  9  1  0 10 11  1  6],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -2741.  -2620.  32184.   1847. -19482.  -7447.  37532. -21924.], 
        // Q{mac}=[ 0  0 31  1  0  0 36  0]

        sign=8'b10011001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00001001, 8'b00000001, 8'b00000000, 8'b00001010, 8'b00001011, 8'b00000001, 8'b00000110};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 141: 
        // x=-117, 
        // s=[-1. -1.  1. -1. -1. -1.  1.  1.],
        // w=[14  2  5 13  2  2  1  6],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -1103.  -2386.  31599.   3368. -19248.  -7213.  37415. -22626.], 
        // Q{mac}=[ 0  0 30  3  0  0 36  0]

        sign=8'b00100011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001110, 8'b00000010, 8'b00000101, 8'b00001101, 8'b00000010, 8'b00000010, 8'b00000001, 8'b00000110};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001011;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 142: 
        // x=-123, 
        // s=[-1.  1.  1. -1. -1.  1. -1. -1.],
        // w=[ 1  0  3 17  7 22  3  1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  -980.  -2386.  31230.   5459. -18387.  -9919.  37784. -22503.], 
        // Q{mac}=[ 0  0 30  5  0  0 36  0]

        sign=8'b01100100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00000000, 8'b00000011, 8'b00010001, 8'b00000111, 8'b00010110, 8'b00000011, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 143: 
        // x=98, 
        // s=[-1. -1. -1.  1.  1. -1.  1. -1.],
        // w=[27 28 42 30 26 37 55  1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -3626.  -5130.  27114.   8399. -15839. -13545.  43174. -22601.], 
        // Q{mac}=[ 0  0 26  8  0  0 42  0]

        sign=8'b00011010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00011011, 8'b00011100, 8'b00101010, 8'b00011110, 8'b00011010, 8'b00100101, 8'b00110111, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b01100010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 144: 
        // x=-35, 
        // s=[ 1.  1. -1. -1. -1. -1. -1.  1.],
        // w=[18 13 13 29 15  6  4  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -4256.  -5585.  27569.   9414. -15314. -13335.  43314. -22706.], 
        // Q{mac}=[ 0  0 26  9  0  0 42  0]

        sign=8'b11000001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00010010, 8'b00001101, 8'b00001101, 8'b00011101, 8'b00001111, 8'b00000110, 8'b00000100, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11011101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 145: 
        // x=57, 
        // s=[ 1.  1.  1. -1.  1.  1. -1.  1.],
        // w=[ 9 13 15 15 20 11 13  0],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -3743.  -4844.  28424.   8559. -14174. -12708.  42573. -22706.], 
        // Q{mac}=[ 0  0 27  8  0  0 41  0]

        sign=8'b11101101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001001, 8'b00001101, 8'b00001111, 8'b00001111, 8'b00010100, 8'b00001011, 8'b00001101, 8'b00000000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00111001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 146: 
        // x=-11, 
        // s=[ 1.  1.  1. -1. -1.  1. -1. -1.],
        // w=[37 36 36 12 17  8 74  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -4150.  -5240.  28028.   8691. -13987. -12796.  43387. -22651.], 
        // Q{mac}=[ 0  0 27  8  0  0 42  0]

        sign=8'b11100100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00100101, 8'b00100100, 8'b00100100, 8'b00001100, 8'b00010001, 8'b00001000, 8'b01001010, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11110101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 147: 
        // x=-3, 
        // s=[-1. -1. -1. -1.  1.  1.  1. -1.],
        // w=[ 2  4 12 14  3  6 20  6],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -4144.  -5228.  28064.   8733. -13996. -12814.  43327. -22633.], 
        // Q{mac}=[ 0  0 27  8  0  0 42  0]

        sign=8'b00001110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00000100, 8'b00001100, 8'b00001110, 8'b00000011, 8'b00000110, 8'b00010100, 8'b00000110};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11111101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 148: 
        // x=29, 
        // s=[-1. -1. -1.  1.  1. -1.  1. -1.],
        // w=[29 29  3 12  7 16 23  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -4985.  -6069.  27977.   9081. -13793. -13278.  43994. -22691.], 
        // Q{mac}=[ 0  0 27  8  0  0 42  0]

        sign=8'b00011010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00011101, 8'b00011101, 8'b00000011, 8'b00001100, 8'b00000111, 8'b00010000, 8'b00010111, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00011101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 149: 
        // x=-26, 
        // s=[-1. -1. -1.  1.  1. -1.  1. -1.],
        // w=[12 22  2 15 15 12  7  9],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -4673.  -5497.  28029.   8691. -14183. -12966.  43812. -22457.], 
        // Q{mac}=[ 0  0 27  8  0  0 42  0]

        sign=8'b00011010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001100, 8'b00010110, 8'b00000010, 8'b00001111, 8'b00001111, 8'b00001100, 8'b00000111, 8'b00001001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11100110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 150: 
        // x=3, 
        // s=[-1. -1. -1. -1. -1. -1.  1.  1.],
        // w=[12 28 30  4 10 10 43  8],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -4709.  -5581.  27939.   8679. -14213. -12996.  43941. -22433.], 
        // Q{mac}=[ 0  0 27  8  0  0 42  0]

        sign=8'b00000011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001100, 8'b00011100, 8'b00011110, 8'b00000100, 8'b00001010, 8'b00001010, 8'b00101011, 8'b00001000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00000011;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 151: 
        // x=-11, 
        // s=[ 1.  1.  1.  1.  1.  1. -1. -1.],
        // w=[15 20 24  6  4 15 28  7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -4874.  -5801.  27675.   8613. -14257. -13161.  44249. -22356.], 
        // Q{mac}=[ 0  0 27  8  0  0 43  0]

        sign=8'b11111100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001111, 8'b00010100, 8'b00011000, 8'b00000110, 8'b00000100, 8'b00001111, 8'b00011100, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11110101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 152: 
        // x=30, 
        // s=[-1. -1. -1.  1.  1. -1.  1. -1.],
        // w=[16 20 12 12 37 37 30  4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -5354.  -6401.  27315.   8973. -13147. -14271.  45149. -22476.], 
        // Q{mac}=[ 0  0 26  8  0  0 44  0]

        sign=8'b00011010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00010000, 8'b00010100, 8'b00001100, 8'b00001100, 8'b00100101, 8'b00100101, 8'b00011110, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00011110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 153: 
        // x=27, 
        // s=[ 1. -1.  1.  1. -1. -1.  1.  1.],
        // w=[1 7 5 9 5 9 3 3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -5327.  -6590.  27450.   9216. -13282. -14514.  45230. -22395.], 
        // Q{mac}=[ 0  0 26  9  0  0 44  0]

        sign=8'b10110011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00000111, 8'b00000101, 8'b00001001, 8'b00000101, 8'b00001001, 8'b00000011, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00011011;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 154: 
        // x=-37, 
        // s=[ 1.  1. -1. -1.  1.  1. -1.  1.],
        // w=[ 1 13  2 14  5 22  9  6],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -5364.  -7071.  27524.   9734. -13467. -15328.  45563. -22617.], 
        // Q{mac}=[ 0  0 26  9  0  0 44  0]

        sign=8'b11001101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00001101, 8'b00000010, 8'b00001110, 8'b00000101, 8'b00010110, 8'b00001001, 8'b00000110};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11011011;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 155: 
        // x=31, 
        // s=[-1. -1. -1.  1. -1. -1.  1.  1.],
        // w=[ 6  6 11  1  1 20 18  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -5550.  -7257.  27183.   9765. -13498. -15948.  46121. -22524.], 
        // Q{mac}=[ 0  0 26  9  0  0 45  0]

        sign=8'b00010011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000110, 8'b00000110, 8'b00001011, 8'b00000001, 8'b00000001, 8'b00010100, 8'b00010010, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00011111;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 156: 
        // x=1, 
        // s=[-1. -1.  1.  1.  1. -1.  1. -1.],
        // w=[ 3 28  5 50 35 34 12  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -5553.  -7285.  27188.   9815. -13463. -15982.  46133. -22529.], 
        // Q{mac}=[ 0  0 26  9  0  0 45  0]

        sign=8'b00111010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00011100, 8'b00000101, 8'b00110010, 8'b00100011, 8'b00100010, 8'b00001100, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00000001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 157: 
        // x=82, 
        // s=[ 1. -1.  1. -1. -1.  1.  1.  1.],
        // w=[ 0 10  9 11 35 15  6  1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -5553.  -8105.  27926.   8913. -16333. -14752.  46625. -22447.], 
        // Q{mac}=[ 0  0 27  8  0  0 45  0]

        sign=8'b10100111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000000, 8'b00001010, 8'b00001001, 8'b00001011, 8'b00100011, 8'b00001111, 8'b00000110, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b01010010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 158: 
        // x=-31, 
        // s=[ 1.  1. -1. -1.  1. -1. -1.  1.],
        // w=[12 24  8  8 36 12 28  0],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -5925.  -8849.  28174.   9161. -17449. -14380.  47493. -22447.], 
        // Q{mac}=[ 0  0 27  8  0  0 46  0]

        sign=8'b11001001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001100, 8'b00011000, 8'b00001000, 8'b00001000, 8'b00100100, 8'b00001100, 8'b00011100, 8'b00000000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11100001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 159: 
        // x=-39, 
        // s=[ 1. -1.  1.  1. -1.  1. -1. -1.],
        // w=[ 6 22  0 41  7 15  2  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -6159.  -7991.  28174.   7562. -17176. -14965.  47571. -22252.], 
        // Q{mac}=[ 0  0 27  7  0  0 46  0]

        sign=8'b10110100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000110, 8'b00010110, 8'b00000000, 8'b00101001, 8'b00000111, 8'b00001111, 8'b00000010, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11011001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 160: 
        // x=-27, 
        // s=[ 1.  1.  1. -1. -1. -1.  1.  1.],
        // w=[ 6  4  1  9 10  2  1  8],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -6321.  -8099.  28147.   7805. -16906. -14911.  47544. -22468.], 
        // Q{mac}=[ 0  0 27  7  0  0 46  0]

        sign=8'b11100011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000110, 8'b00000100, 8'b00000001, 8'b00001001, 8'b00001010, 8'b00000010, 8'b00000001, 8'b00001000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11100101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 161: 
        // x=-23, 
        // s=[-1.  1.  1.  1.  1. -1. -1.  1.],
        // w=[15  6  4 13  9 14  3  8],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -5976.  -8237.  28055.   7506. -17113. -14589.  47613. -22652.], 
        // Q{mac}=[ 0  0 27  7  0  0 46  0]

        sign=8'b01111001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001111, 8'b00000110, 8'b00000100, 8'b00001101, 8'b00001001, 8'b00001110, 8'b00000011, 8'b00001000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11101001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 162: 
        // x=-13, 
        // s=[-1. -1. -1.  1.  1. -1. -1.  1.],
        // w=[ 2  4 11 11  6 14  1  8],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -5950.  -8185.  28198.   7363. -17191. -14407.  47626. -22756.], 
        // Q{mac}=[ 0  0 27  7  0  0 46  0]

        sign=8'b00011001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00000100, 8'b00001011, 8'b00001011, 8'b00000110, 8'b00001110, 8'b00000001, 8'b00001000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11110011;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 163: 
        // x=-116, 
        // s=[ 1. -1.  1.  1. -1. -1.  1.  1.],
        // w=[ 0 13 14  4  5  2  6  1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -5950.  -6677.  26574.   6899. -16611. -14175.  46930. -22872.], 
        // Q{mac}=[ 0  0 25  6  0  0 45  0]

        sign=8'b10110011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000000, 8'b00001101, 8'b00001110, 8'b00000100, 8'b00000101, 8'b00000010, 8'b00000110, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001100;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 164: 
        // x=-117, 
        // s=[-1.  1. -1.  1.  1.  1. -1.  1.],
        // w=[7 2 3 6 1 5 9 8],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -5131.  -6911.  26925.   6197. -16728. -14760.  47983. -23808.], 
        // Q{mac}=[ 0  0 26  6  0  0 46  0]

        sign=8'b01011101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00000010, 8'b00000011, 8'b00000110, 8'b00000001, 8'b00000101, 8'b00001001, 8'b00001000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001011;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 165: 
        // x=-121, 
        // s=[ 1. -1.  1. -1.  1. -1. -1.  1.],
        // w=[ 0  6  5  3 12  3  2  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -5131.  -6185.  26320.   6560. -18180. -14397.  48225. -24050.], 
        // Q{mac}=[ 0  0 25  6  0  0 47  0]

        sign=8'b10101001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000000, 8'b00000110, 8'b00000101, 8'b00000011, 8'b00001100, 8'b00000011, 8'b00000010, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000111;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 166: 
        // x=-117, 
        // s=[-1. -1.  1. -1.  1.  1.  1. -1.],
        // w=[14 14 13  1  1  3  5  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -3493.  -4547.  24799.   6677. -18297. -14748.  47640. -23816.], 
        // Q{mac}=[ 0  0 24  6  0  0 46  0]

        sign=8'b00101110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001110, 8'b00001110, 8'b00001101, 8'b00000001, 8'b00000001, 8'b00000011, 8'b00000101, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001011;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 167: 
        // x=-119, 
        // s=[-1.  1.  1.  1.  1.  1. -1.  1.],
        // w=[4 4 2 2 6 4 7 3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -3017.  -5023.  24561.   6439. -19011. -15224.  48473. -24173.], 
        // Q{mac}=[ 0  0 23  6  0  0 47  0]

        sign=8'b01111101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000100, 8'b00000100, 8'b00000010, 8'b00000010, 8'b00000110, 8'b00000100, 8'b00000111, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 168: 
        // x=-123, 
        // s=[-1.  1.  1. -1.  1. -1. -1. -1.],
        // w=[ 4  4  3  1 11  3  3  1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -2525.  -5515.  24192.   6562. -20364. -14855.  48842. -24050.], 
        // Q{mac}=[ 0  0 23  6  0  0 47  0]

        sign=8'b01101000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000100, 8'b00000100, 8'b00000011, 8'b00000001, 8'b00001011, 8'b00000011, 8'b00000011, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 169: 
        // x=-112, 
        // s=[ 1. -1.  1. -1. -1.  1.  1.  1.],
        // w=[ 2 13  2  7 15 10  7  9],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -2749.  -4059.  23968.   7346. -18684. -15975.  48058. -25058.], 
        // Q{mac}=[ 0  0 23  7  0  0 46  0]

        sign=8'b10100111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00001101, 8'b00000010, 8'b00000111, 8'b00001111, 8'b00001010, 8'b00000111, 8'b00001001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10010000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 170: 
        // x=-117, 
        // s=[-1.  1.  1. -1.  1.  1. -1. -1.],
        // w=[11  2  2  2  4  1  8  4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -1462.  -4293.  23734.   7580. -19152. -16092.  48994. -24590.], 
        // Q{mac}=[ 0  0 23  7  0  0 47  0]

        sign=8'b01101100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001011, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000100, 8'b00000001, 8'b00001000, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001011;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 171: 
        // x=-115, 
        // s=[-1.  1. -1. -1.  1. -1.  1. -1.],
        // w=[ 2  8  3  7 18  4  5  4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ -1232.  -5213.  24079.   8385. -21222. -15632.  48419. -24130.], 
        // Q{mac}=[ 0  0 23  8  0  0 47  0]

        sign=8'b01001010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00001000, 8'b00000011, 8'b00000111, 8'b00010010, 8'b00000100, 8'b00000101, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 172: 
        // x=114, 
        // s=[ 1.  1.  1.  1.  1. -1.  1.  1.],
        // w=[ 5 15  0  5  5  4  2  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  -662.  -3503.  24079.   8955. -20652. -16088.  48647. -23788.], 
        // Q{mac}=[ 0  0 23  8  0  0 47  0]

        sign=8'b11111011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000101, 8'b00001111, 8'b00000000, 8'b00000101, 8'b00000101, 8'b00000100, 8'b00000010, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b01110010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 173: 
        // x=116, 
        // s=[ 1. -1.  1.  1.  1.  1. -1. -1.],
        // w=[12  5  9 10  6  4  1  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[   730.  -4083.  25123.  10115. -19956. -15624.  48531. -24020.], 
        // Q{mac}=[ 0  0 24  9  0  0 47  0]

        sign=8'b10111100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001100, 8'b00000101, 8'b00001001, 8'b00001010, 8'b00000110, 8'b00000100, 8'b00000001, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b01110100;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 174: 
        // x=120, 
        // s=[-1.  1.  1.  1.  1.  1. -1. -1.],
        // w=[3 1 1 5 5 1 6 8],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[   370.  -3963.  25243.  10715. -19356. -15504.  47811. -24980.], 
        // Q{mac}=[ 0  0 24 10  0  0 46  0]

        sign=8'b01111100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00000001, 8'b00000001, 8'b00000101, 8'b00000101, 8'b00000001, 8'b00000110, 8'b00001000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b01111000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 175: 
        // x=-120, 
        // s=[-1. -1.  1. -1. -1. -1. -1.  1.],
        // w=[14  1  9  9  6  3  7  1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  2050.  -3843.  24163.  11795. -18636. -15144.  48651. -25100.], 
        // Q{mac}=[ 2  0 23 11  0  0 47  0]

        sign=8'b00100001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001110, 8'b00000001, 8'b00001001, 8'b00001001, 8'b00000110, 8'b00000011, 8'b00000111, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 176: 
        // x=-128, 
        // s=[-1. -1.  1. -1.  1.  1. -1.  1.],
        // w=[7 1 0 6 0 7 9 8],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  2946.  -3715.  24163.  12563. -18636. -16040.  49803. -26124.], 
        // Q{mac}=[ 2  0 23 12  0  0 48  0]

        sign=8'b00101101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00000001, 8'b00000000, 8'b00000110, 8'b00000000, 8'b00000111, 8'b00001001, 8'b00001000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 177: 
        // x=-128, 
        // s=[ 1. -1. -1. -1. -1.  1. -1.  1.],
        // w=[1 7 4 8 2 3 6 9],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  2818.  -2819.  24675.  13587. -18380. -16424.  50571. -27276.], 
        // Q{mac}=[ 2  0 24 13  0  0 49  0]

        sign=8'b10000101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00000111, 8'b00000100, 8'b00001000, 8'b00000010, 8'b00000011, 8'b00000110, 8'b00001001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 178: 
        // x=-128, 
        // s=[-1.  1. -1.  1. -1. -1. -1. -1.],
        // w=[10  0  4  2  5  7  3  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  4098.  -2819.  25187.  13331. -17740. -15528.  50955. -26636.], 
        // Q{mac}=[ 4  0 24 13  0  0 49  0]

        sign=8'b01010000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001010, 8'b00000000, 8'b00000100, 8'b00000010, 8'b00000101, 8'b00000111, 8'b00000011, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 179: 
        // x=-120, 
        // s=[-1. -1.  1.  1. -1. -1.  1. -1.],
        // w=[11 15 14  1  8  3  7  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  5418.  -1019.  23507.  13211. -16780. -15168.  50115. -26396.], 
        // Q{mac}=[ 5  0 22 12  0  0 48  0]

        sign=8'b00110010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001011, 8'b00001111, 8'b00001110, 8'b00000001, 8'b00001000, 8'b00000011, 8'b00000111, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 180: 
        // x=-123, 
        // s=[-1.  1. -1.  1.  1. -1.  1.  1.],
        // w=[2 4 8 1 8 2 0 1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  5664.  -1511.  24491.  13088. -17764. -14922.  50115. -26519.], 
        // Q{mac}=[ 5  0 23 12  0  0 48  0]

        sign=8'b01011011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00000100, 8'b00001000, 8'b00000001, 8'b00001000, 8'b00000010, 8'b00000000, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 181: 
        // x=-125, 
        // s=[-1.  1. -1.  1.  1. -1. -1. -1.],
        // w=[ 7  2  1  2 14 13  5  4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  6539.  -1761.  24616.  12838. -19514. -13297.  50740. -26019.], 
        // Q{mac}=[ 6  0 24 12  0  0 49  0]

        sign=8'b01011000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00000010, 8'b00000001, 8'b00000010, 8'b00001110, 8'b00001101, 8'b00000101, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000011;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 182: 
        // x=4, 
        // s=[-1. -1. -1.  1.  1. -1.  1. -1.],
        // w=[41 40 22 15 21 15 54  6],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  6375.  -1921.  24528.  12898. -19430. -13357.  50956. -26043.], 
        // Q{mac}=[ 6  0 23 12  0  0 49  0]

        sign=8'b00011010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00101001, 8'b00101000, 8'b00010110, 8'b00001111, 8'b00010101, 8'b00001111, 8'b00110110, 8'b00000110};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00000100;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 183: 
        // x=9, 
        // s=[-1.  1. -1. -1.  1.  1. -1.  1.],
        // w=[ 2 30  1 11 10  0 16  0],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  6357.  -1651.  24519.  12799. -19340. -13357.  50812. -26043.], 
        // Q{mac}=[ 6  0 23 12  0  0 49  0]

        sign=8'b01001101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00011110, 8'b00000001, 8'b00001011, 8'b00001010, 8'b00000000, 8'b00010000, 8'b00000000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00001001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 184: 
        // x=-26, 
        // s=[-1. -1.  1. -1. -1.  1.  1. -1.],
        // w=[18  6  3  4  5  8  1  6],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  6825.  -1495.  24441.  12903. -19210. -13565.  50786. -25887.], 
        // Q{mac}=[ 6  0 23 12  0  0 49  0]

        sign=8'b00100110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00010010, 8'b00000110, 8'b00000011, 8'b00000100, 8'b00000101, 8'b00001000, 8'b00000001, 8'b00000110};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11100110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 185: 
        // x=13, 
        // s=[ 1.  1.  1. -1. -1.  1. -1. -1.],
        // w=[48 58 30 23 14 28 94  4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  7449.   -741.  24831.  12604. -19392. -13201.  49564. -25939.], 
        // Q{mac}=[ 7  0 24 12  0  0 48  0]

        sign=8'b11100100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00110000, 8'b00111010, 8'b00011110, 8'b00010111, 8'b00001110, 8'b00011100, 8'b01011110, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00001101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 186: 
        // x=-4, 
        // s=[ 1.  1.  1. -1. -1.  1. -1. -1.],
        // w=[50 69  8 41 11 44 75  1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  7249.  -1017.  24799.  12768. -19348. -13377.  49864. -25935.], 
        // Q{mac}=[ 7  0 24 12  0  0 48  0]

        sign=8'b11100100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00110010, 8'b01000101, 8'b00001000, 8'b00101001, 8'b00001011, 8'b00101100, 8'b01001011, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11111100;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 187: 
        // x=24, 
        // s=[ 1.  1.  1. -1. -1.  1. -1. -1.],
        // w=[37 43 34 18 10 24 47  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 8.1370e+03  1.5000e+01  2.5615e+04  1.2336e+04 -1.9588e+04 -1.2801e+04    4.8736e+04 -2.6055e+04], 
        // Q{mac}=[ 7  0 25 12  0  0 47  0]

        sign=8'b11100100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00100101, 8'b00101011, 8'b00100010, 8'b00010010, 8'b00001010, 8'b00011000, 8'b00101111, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00011000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 188: 
        // x=38, 
        // s=[-1.  1.  1.  1. -1. -1.  1.  1.],
        // w=[21  2  4  5  1  6  8  0],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  7339.     91.  25767.  12526. -19626. -13029.  49040. -26055.], 
        // Q{mac}=[ 7  0 25 12  0  0 47  0]

        sign=8'b01110011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00010101, 8'b00000010, 8'b00000100, 8'b00000101, 8'b00000001, 8'b00000110, 8'b00001000, 8'b00000000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00100110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 189: 
        // x=14, 
        // s=[-1. -1. -1. -1. -1. -1.  1. -1.],
        // w=[ 5 20 35  6 14  8 54  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  7269.   -189.  25277.  12442. -19822. -13141.  49796. -26083.], 
        // Q{mac}=[ 7  0 24 12  0  0 48  0]

        sign=8'b00000010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000101, 8'b00010100, 8'b00100011, 8'b00000110, 8'b00001110, 8'b00001000, 8'b00110110, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00001110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 190: 
        // x=6, 
        // s=[ 1. -1. -1.  1. -1.  1.  1. -1.],
        // w=[ 5 17 14 16 27 17  3  4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  7299.   -291.  25193.  12538. -19984. -13039.  49814. -26107.], 
        // Q{mac}=[ 7  0 24 12  0  0 48  0]

        sign=8'b10010110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000101, 8'b00010001, 8'b00001110, 8'b00010000, 8'b00011011, 8'b00010001, 8'b00000011, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00000110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 191: 
        // x=8, 
        // s=[ 1.  1. -1.  1.  1.  1.  1. -1.],
        // w=[ 7 11  5  3  4  3  1  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  7355.   -203.  25153.  12562. -19952. -13015.  49822. -26123.], 
        // Q{mac}=[ 7  0 24 12  0  0 48  0]

        sign=8'b11011110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00001011, 8'b00000101, 8'b00000011, 8'b00000100, 8'b00000011, 8'b00000001, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00001000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 192: 
        // x=24, 
        // s=[-1. -1. -1.  1. -1.  1.  1.  1.],
        // w=[27 55 22 23 27 12 56  4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  6707.  -1523.  24625.  13114. -20600. -12727.  51166. -26027.], 
        // Q{mac}=[ 6  0 24 12  0  0 49  0]

        sign=8'b00010111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00011011, 8'b00110111, 8'b00010110, 8'b00010111, 8'b00011011, 8'b00001100, 8'b00111000, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00011000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 193: 
        // x=39, 
        // s=[ 1. -1. -1. -1. -1.  1.  1. -1.],
        // w=[18  8  5  8 28 18  6  1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  7409.  -1835.  24430.  12802. -21692. -12025.  51400. -26066.], 
        // Q{mac}=[ 7  0 23 12  0  0 50  0]

        sign=8'b10000110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00010010, 8'b00001000, 8'b00000101, 8'b00001000, 8'b00011100, 8'b00010010, 8'b00000110, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00100111;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 194: 
        // x=-28, 
        // s=[ 1.  1. -1. -1. -1.  1. -1.  1.],
        // w=[15 18  7 10 13 45 14  4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  6989.  -2339.  24626.  13082. -21328. -13285.  51792. -26178.], 
        // Q{mac}=[ 6  0 24 12  0  0 50  0]

        sign=8'b11000101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001111, 8'b00010010, 8'b00000111, 8'b00001010, 8'b00001101, 8'b00101101, 8'b00001110, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11100100;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 195: 
        // x=21, 
        // s=[ 1.  1. -1. -1. -1.  1. -1.  1.],
        // w=[ 7 16  7 24 13  5  2  1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  7136.  -2003.  24479.  12578. -21601. -13180.  51750. -26157.], 
        // Q{mac}=[ 6  0 23 12  0  0 50  0]

        sign=8'b11000101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00010000, 8'b00000111, 8'b00011000, 8'b00001101, 8'b00000101, 8'b00000010, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00010101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 196: 
        // x=18, 
        // s=[-1. -1. -1.  1. -1. -1.  1.  1.],
        // w=[21 29  9 21  4 18 29  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  6758.  -2525.  24317.  12956. -21673. -13504.  52272. -26121.], 
        // Q{mac}=[ 6  0 23 12  0  0 51  0]

        sign=8'b00010011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00010101, 8'b00011101, 8'b00001001, 8'b00010101, 8'b00000100, 8'b00010010, 8'b00011101, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00010010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 197: 
        // x=15, 
        // s=[ 1.  1. -1.  1.  1. -1. -1. -1.],
        // w=[10 46 13  7 58 42 33 12],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  6908.  -1835.  24122.  13061. -20803. -14134.  51777. -26301.], 
        // Q{mac}=[ 6  0 23 12  0  0 50  0]

        sign=8'b11011000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001010, 8'b00101110, 8'b00001101, 8'b00000111, 8'b00111010, 8'b00101010, 8'b00100001, 8'b00001100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00001111;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 198: 
        // x=-21, 
        // s=[-1. -1.  1.  1.  1. -1. -1. -1.],
        // w=[18 11 30 35 80 61 35  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  7286.  -1604.  23492.  12326. -22483. -12853.  52512. -26259.], 
        // Q{mac}=[ 7  0 22 12  0  0 51  0]

        sign=8'b00111000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00010010, 8'b00001011, 8'b00011110, 8'b00100011, 8'b01010000, 8'b00111101, 8'b00100011, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11101011;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 199: 
        // x=-42, 
        // s=[-1. -1.  1.  1.  1. -1. -1. -1.],
        // w=[26  8 33 13 40 33 22  8],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  8378.  -1268.  22106.  11780. -24163. -11467.  53436. -25923.], 
        // Q{mac}=[ 8  0 21 11  0  0 52  0]

        sign=8'b00111000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00011010, 8'b00001000, 8'b00100001, 8'b00001101, 8'b00101000, 8'b00100001, 8'b00010110, 8'b00001000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11010110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 200: 
        // x=-112, 
        // s=[-1.  1.  1. -1. -1.  1.  1.  1.],
        // w=[11  1  2  2  1 18  3  6],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  9610.  -1380.  21882.  12004. -24051. -13483.  53100. -26595.], 
        // Q{mac}=[ 9  0 21 11  0  0 51  0]

        sign=8'b01100111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001011, 8'b00000001, 8'b00000010, 8'b00000010, 8'b00000001, 8'b00010010, 8'b00000011, 8'b00000110};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10010000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 201: 
        // x=-91, 
        // s=[ 1.  1. -1. -1.  1.  1.  1.  1.],
        // w=[10 12 14 10  1  6  4 11],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  8700.  -2472.  23156.  12914. -24142. -14029.  52736. -27596.], 
        // Q{mac}=[ 8  0 22 12  0  0 51  0]

        sign=8'b11001111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001010, 8'b00001100, 8'b00001110, 8'b00001010, 8'b00000001, 8'b00000110, 8'b00000100, 8'b00001011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10100101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 202: 
        // x=-96, 
        // s=[ 1.  1. -1. -1.  1.  1.  1.  1.],
        // w=[13 18 15  7  1  6  4  1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  7452.  -4200.  24596.  13586. -24238. -14605.  52352. -27692.], 
        // Q{mac}=[ 7  0 24 13  0  0 51  0]

        sign=8'b11001111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001101, 8'b00010010, 8'b00001111, 8'b00000111, 8'b00000001, 8'b00000110, 8'b00000100, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10100000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 203: 
        // x=-98, 
        // s=[ 1.  1. -1. -1.  1.  1.  1.  1.],
        // w=[ 7 12 20 10 11  7  7  1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  6766.  -5376.  26556.  14566. -25316. -15291.  51666. -27790.], 
        // Q{mac}=[ 6  0 25 14  0  0 50  0]

        sign=8'b11001111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00001100, 8'b00010100, 8'b00001010, 8'b00001011, 8'b00000111, 8'b00000111, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10011110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 204: 
        // x=-126, 
        // s=[-1.  1.  1. -1.  1. -1.  1.  1.],
        // w=[7 0 8 9 8 2 3 5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  7648.  -5376.  25548.  15700. -26324. -15039.  51288. -28420.], 
        // Q{mac}=[ 7  0 24 15  0  0 50  0]

        sign=8'b01101011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00000000, 8'b00001000, 8'b00001001, 8'b00001000, 8'b00000010, 8'b00000011, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 205: 
        // x=-112, 
        // s=[-1.  1. -1.  1. -1.  1. -1. -1.],
        // w=[8 8 9 0 6 4 2 3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  8544.  -6272.  26556.  15700. -25652. -15487.  51512. -28084.], 
        // Q{mac}=[ 8  0 25 15  0  0 50  0]

        sign=8'b01010100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001000, 8'b00001000, 8'b00001001, 8'b00000000, 8'b00000110, 8'b00000100, 8'b00000010, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10010000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 206: 
        // x=-126, 
        // s=[-1.  1. -1. -1. -1. -1. -1.  1.],
        // w=[4 6 7 3 6 5 3 9],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  9048.  -7028.  27438.  16078. -24896. -14857.  51890. -29218.], 
        // Q{mac}=[ 8  0 26 15  0  0 50  0]

        sign=8'b01000001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000100, 8'b00000110, 8'b00000111, 8'b00000011, 8'b00000110, 8'b00000101, 8'b00000011, 8'b00001001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 207: 
        // x=-111, 
        // s=[ 1.  1. -1.  1. -1.  1. -1.  1.],
        // w=[ 0 10  1  4 10  4  2  1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  9048.  -8138.  27549.  15634. -23786. -15301.  52112. -29329.], 
        // Q{mac}=[ 8  0 26 15  0  0 50  0]

        sign=8'b11010101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000000, 8'b00001010, 8'b00000001, 8'b00000100, 8'b00001010, 8'b00000100, 8'b00000010, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10010001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 208: 
        // x=32, 
        // s=[-1.  1. -1.  1.  1.  1. -1. -1.],
        // w=[1 6 6 4 2 0 9 3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  9016.  -7946.  27357.  15762. -23722. -15301.  51824. -29425.], 
        // Q{mac}=[ 8  0 26 15  0  0 50  0]

        sign=8'b01011100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00000110, 8'b00000110, 8'b00000100, 8'b00000010, 8'b00000000, 8'b00001001, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00100000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 209: 
        // x=6, 
        // s=[-1. -1.  1.  1.  1. -1. -1.  1.],
        // w=[16 17  8 15 12 15  5  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  8920.  -8048.  27405.  15852. -23650. -15391.  51794. -29413.], 
        // Q{mac}=[ 8  0 26 15  0  0 50  0]

        sign=8'b00111001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00010000, 8'b00010001, 8'b00001000, 8'b00001111, 8'b00001100, 8'b00001111, 8'b00000101, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00000110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 210: 
        // x=-27, 
        // s=[ 1.  1. -1. -1. -1.  1.  1.  1.],
        // w=[18 10  8 12  1  1 13  0],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  8434.  -8318.  27621.  16176. -23623. -15418.  51443. -29413.], 
        // Q{mac}=[ 8  0 26 15  0  0 50  0]

        sign=8'b11000111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00010010, 8'b00001010, 8'b00001000, 8'b00001100, 8'b00000001, 8'b00000001, 8'b00001101, 8'b00000000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11100101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 211: 
        // x=77, 
        // s=[ 1.  1. -1. -1. -1.  1.  1. -1.],
        // w=[ 1 14  1 13  1 11  8  8],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  8511.  -7240.  27544.  15175. -23700. -14571.  52059. -30029.], 
        // Q{mac}=[ 8  0 26 14  0  0 50  0]

        sign=8'b11000110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00001110, 8'b00000001, 8'b00001101, 8'b00000001, 8'b00001011, 8'b00001000, 8'b00001000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b01001101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 212: 
        // x=-73, 
        // s=[ 1.  1.  1. -1. -1.  1. -1.  1.],
        // w=[ 4 12  1 14 14  9  1  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  8219.  -8116.  27471.  16197. -22678. -15228.  52132. -30248.], 
        // Q{mac}=[ 8  0 26 15  0  0 50  0]

        sign=8'b11100101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000100, 8'b00001100, 8'b00000001, 8'b00001110, 8'b00001110, 8'b00001001, 8'b00000001, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10110111;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 213: 
        // x=-112, 
        // s=[-1. -1. -1.  1. -1.  1.  1.  1.],
        // w=[11  5  7  0  4  5 13  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  9451.  -7556.  28255.  16197. -22230. -15788.  50676. -30584.], 
        // Q{mac}=[ 9  0 27 15  0  0 49  0]

        sign=8'b00010111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001011, 8'b00000101, 8'b00000111, 8'b00000000, 8'b00000100, 8'b00000101, 8'b00001101, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10010000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 214: 
        // x=-91, 
        // s=[ 1.  1. -1. -1.  1.  1.  1.  1.],
        // w=[ 2 12 13  8  7  0  1 12],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  9269.  -8648.  29438.  16925. -22867. -15788.  50585. -31676.], 
        // Q{mac}=[ 9  0 28 16  0  0 49  0]

        sign=8'b11001111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00001100, 8'b00001101, 8'b00001000, 8'b00000111, 8'b00000000, 8'b00000001, 8'b00001100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10100101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 215: 
        // x=-96, 
        // s=[-1.  1. -1.  1. -1. -1. -1.  1.],
        // w=[ 1  8 15  0  1  3  3  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  9365.  -9416.  30878.  16925. -22771. -15500.  50873. -31868.], 
        // Q{mac}=[ 9  0 30 16  0  0 49  0]

        sign=8'b01010001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00001000, 8'b00001111, 8'b00000000, 8'b00000001, 8'b00000011, 8'b00000011, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10100000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 216: 
        // x=-98, 
        // s=[ 1.  1. -1. -1.  1.  1.  1.  1.],
        // w=[ 6 10 17 12 11  8  7  8],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  8777. -10396.  32544.  18101. -23849. -16284.  50187. -32652.], 
        // Q{mac}=[ 8  0 31 17  0  0 49  0]

        sign=8'b11001111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000110, 8'b00001010, 8'b00010001, 8'b00001100, 8'b00001011, 8'b00001000, 8'b00000111, 8'b00001000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10011110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 217: 
        // x=-126, 
        // s=[-1. -1.  1.  1. -1. -1. -1.  1.],
        // w=[1 5 1 1 3 8 3 4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  8903.  -9766.  32418.  17975. -23471. -15276.  50565. -33156.], 
        // Q{mac}=[ 8  0 31 17  0  0 49  0]

        sign=8'b00110001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00000101, 8'b00000001, 8'b00000001, 8'b00000011, 8'b00001000, 8'b00000011, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 218: 
        // x=-112, 
        // s=[-1.  1.  1. -1. -1.  1.  1.  1.],
        // w=[ 6  7  0  5  6 17  6  7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  9575. -10550.  32418.  18535. -22799. -17180.  49893. -33940.], 
        // Q{mac}=[ 9  0 31 18  0  0 48  0]

        sign=8'b01100111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000110, 8'b00000111, 8'b00000000, 8'b00000101, 8'b00000110, 8'b00010001, 8'b00000110, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10010000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 219: 
        // x=-126, 
        // s=[ 1.  1. -1. -1. -1. -1. -1. -1.],
        // w=[ 7  6  6 11  4  1  1  1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  8693. -11306.  33174.  19921. -22295. -17054.  50019. -33814.], 
        // Q{mac}=[ 8  0 32 19  0  0 48  0]

        sign=8'b11000000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00000110, 8'b00000110, 8'b00001011, 8'b00000100, 8'b00000001, 8'b00000001, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 220: 
        // x=-111, 
        // s=[ 1. -1.  1.  1.  1.  1.  1.  1.],
        // w=[1 4 0 8 1 6 1 9],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  8582. -10862.  33174.  19033. -22406. -17720.  49908. -34813.], 
        // Q{mac}=[ 8  0 32 18  0  0 48  0]

        sign=8'b10111111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00000100, 8'b00000000, 8'b00001000, 8'b00000001, 8'b00000110, 8'b00000001, 8'b00001001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10010001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 221: 
        // x=32, 
        // s=[-1.  1. -1. -1.  1.  1. -1.  1.],
        // w=[ 3  3  2  5 12 11  7  7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  8486. -10766.  33110.  18873. -22022. -17368.  49684. -34589.], 
        // Q{mac}=[ 8  0 32 18  0  0 48  0]

        sign=8'b01001101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00000011, 8'b00000010, 8'b00000101, 8'b00001100, 8'b00001011, 8'b00000111, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00100000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 222: 
        // x=6, 
        // s=[-1. -1.  1.  1.  1. -1. -1.  1.],
        // w=[22 14  9 16  5 15 13  9],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  8354. -10850.  33164.  18969. -21992. -17458.  49606. -34535.], 
        // Q{mac}=[ 8  0 32 18  0  0 48  0]

        sign=8'b00111001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00010110, 8'b00001110, 8'b00001001, 8'b00010000, 8'b00000101, 8'b00001111, 8'b00001101, 8'b00001001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00000110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 223: 
        // x=-27, 
        // s=[ 1.  1. -1. -1. -1.  1.  1. -1.],
        // w=[11  0  6  1  5 12  6  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  8057. -10850.  33326.  18996. -21857. -17782.  49444. -34454.], 
        // Q{mac}=[ 7  0 32 18  0  0 48  0]

        sign=8'b11000110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001011, 8'b00000000, 8'b00000110, 8'b00000001, 8'b00000101, 8'b00001100, 8'b00000110, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11100101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 224: 
        // x=77, 
        // s=[-1.  1. -1. -1.  1.  1. -1. -1.],
        // w=[ 3  3 10  6  4 23  3 10],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  7826. -10619.  32556.  18534. -21549. -16011.  49213. -35224.], 
        // Q{mac}=[ 7  0 31 18  0  0 48  0]

        sign=8'b01001100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00000011, 8'b00001010, 8'b00000110, 8'b00000100, 8'b00010111, 8'b00000011, 8'b00001010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b01001101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 225: 
        // x=-73, 
        // s=[ 1.  1. -1.  1. -1.  1. -1.  1.],
        // w=[ 9  6  7  0 13 10 10  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  7169. -11057.  33067.  18534. -20600. -16741.  49943. -35443.], 
        // Q{mac}=[ 7  0 32 18  0  0 48  0]

        sign=8'b11010101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001001, 8'b00000110, 8'b00000111, 8'b00000000, 8'b00001101, 8'b00001010, 8'b00001010, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10110111;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 226: 
        // x=-120, 
        // s=[-1. -1. -1.  1.  1.  1.  1.  1.],
        // w=[ 9  1  2  3 11  2  7 10],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  8249. -10937.  33307.  18174. -21920. -16981.  49103. -36643.], 
        // Q{mac}=[ 8  0 32 17  0  0 47  0]

        sign=8'b00011111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001001, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00001011, 8'b00000010, 8'b00000111, 8'b00001010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 227: 
        // x=-115, 
        // s=[-1. -1. -1. -1.  1.  1.  1.  1.],
        // w=[ 3  2 12  3  6  3  9  4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  8594. -10707.  34687.  18519. -22610. -17326.  48068. -37103.], 
        // Q{mac}=[ 8  0 33 18  0  0 46  0]

        sign=8'b00001111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00000010, 8'b00001100, 8'b00000011, 8'b00000110, 8'b00000011, 8'b00001001, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 228: 
        // x=-116, 
        // s=[ 1.  1. -1. -1.  1. -1.  1.  1.],
        // w=[ 0  9  7  4 23  8  2 11],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  8594. -11751.  35499.  18983. -25278. -16398.  47836. -38379.], 
        // Q{mac}=[ 8  0 34 18  0  0 46  0]

        sign=8'b11001011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000000, 8'b00001001, 8'b00000111, 8'b00000100, 8'b00010111, 8'b00001000, 8'b00000010, 8'b00001011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001100;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 229: 
        // x=-116, 
        // s=[ 1. -1. -1. -1.  1.  1.  1.  1.],
        // w=[4 2 1 9 3 7 6 5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  8130. -11519.  35615.  20027. -25626. -17210.  47140. -38959.], 
        // Q{mac}=[ 7  0 34 19  0  0 46  0]

        sign=8'b10001111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000100, 8'b00000010, 8'b00000001, 8'b00001001, 8'b00000011, 8'b00000111, 8'b00000110, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001100;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 230: 
        // x=-125, 
        // s=[ 1. -1.  1.  1. -1.  1. -1. -1.],
        // w=[ 2 11  3  5  3 10  5  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  7880. -10144.  35240.  19402. -25251. -18460.  47765. -38709.], 
        // Q{mac}=[ 7  0 34 18  0  0 46  0]

        sign=8'b10110100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00001011, 8'b00000011, 8'b00000101, 8'b00000011, 8'b00001010, 8'b00000101, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000011;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 231: 
        // x=-120, 
        // s=[-1.  1.  1. -1.  1.  1.  1.  1.],
        // w=[ 7  1  3  7 14  5  1  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  8720. -10264.  34880.  20242. -26931. -19060.  47645. -39309.], 
        // Q{mac}=[ 8  0 34 19  0  0 46  0]

        sign=8'b01101111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00000001, 8'b00000011, 8'b00000111, 8'b00001110, 8'b00000101, 8'b00000001, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 232: 
        // x=-128, 
        // s=[ 1.  1.  1. -1.  1. -1. -1.  1.],
        // w=[ 4  6  6  3  1 11  4  0],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  8208. -11032.  34112.  20626. -27059. -17652.  48157. -39309.], 
        // Q{mac}=[ 8  0 33 20  0  0 47  0]

        sign=8'b11101001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000100, 8'b00000110, 8'b00000110, 8'b00000011, 8'b00000001, 8'b00001011, 8'b00000100, 8'b00000000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 233: 
        // x=-118, 
        // s=[-1.  1. -1.  1.  1. -1. -1.  1.],
        // w=[10  4 12  5 12  7  3  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  9388. -11504.  35528.  20036. -28475. -16826.  48511. -39899.], 
        // Q{mac}=[ 9  0 34 19  0  0 47  0]

        sign=8'b01011001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001010, 8'b00000100, 8'b00001100, 8'b00000101, 8'b00001100, 8'b00000111, 8'b00000011, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 234: 
        // x=-18, 
        // s=[-1.  1.  1.  1.  1.  1.  1. -1.],
        // w=[ 4  5  1  0  8 11  7  6],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  9460. -11594.  35510.  20036. -28619. -17024.  48385. -39791.], 
        // Q{mac}=[ 9  0 34 19  0  0 47  0]

        sign=8'b01111110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000100, 8'b00000101, 8'b00000001, 8'b00000000, 8'b00001000, 8'b00001011, 8'b00000111, 8'b00000110};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11101110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 235: 
        // x=29, 
        // s=[ 1. -1. -1. -1. -1. -1.  1.  1.],
        // w=[ 5  3  6  2  3  5 11  0],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  9605. -11681.  35336.  19978. -28706. -17169.  48704. -39791.], 
        // Q{mac}=[ 9  0 34 19  0  0 47  0]

        sign=8'b10000011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000101, 8'b00000011, 8'b00000110, 8'b00000010, 8'b00000011, 8'b00000101, 8'b00001011, 8'b00000000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00011101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 236: 
        // x=-45, 
        // s=[ 1.  1.  1. -1. -1.  1.  1.  1.],
        // w=[ 9  2 13 25 17 18  7  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  9200. -11771.  34751.  21103. -27941. -17979.  48389. -39926.], 
        // Q{mac}=[ 8  0 33 20  0  0 47  0]

        sign=8'b11100111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001001, 8'b00000010, 8'b00001101, 8'b00011001, 8'b00010001, 8'b00010010, 8'b00000111, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11010011;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 237: 
        // x=41, 
        // s=[ 1. -1. -1.  1.  1. -1. -1.  1.],
        // w=[ 2  2 16 22 24 37  6  0],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  9282. -11853.  34095.  22005. -26957. -19496.  48143. -39926.], 
        // Q{mac}=[ 9  0 33 21  0  0 47  0]

        sign=8'b10011001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00000010, 8'b00010000, 8'b00010110, 8'b00011000, 8'b00100101, 8'b00000110, 8'b00000000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00101001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 238: 
        // x=-35, 
        // s=[ 1.  1.  1.  1. -1.  1. -1. -1.],
        // w=[17 13 12  5  7  1 26  6],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  8687. -12308.  33675.  21830. -26712. -19531.  49053. -39716.], 
        // Q{mac}=[ 8  0 32 21  0  0 47  0]

        sign=8'b11110100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00010001, 8'b00001101, 8'b00001100, 8'b00000101, 8'b00000111, 8'b00000001, 8'b00011010, 8'b00000110};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11011101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 239: 
        // x=-102, 
        // s=[-1. -1.  1. -1.  1.  1. -1.  1.],
        // w=[ 9  3  1  5 12  0  1  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  9605. -12002.  33573.  22340. -27936. -19531.  49155. -40226.], 
        // Q{mac}=[ 9  0 32 21  0  0 48  0]

        sign=8'b00101101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001001, 8'b00000011, 8'b00000001, 8'b00000101, 8'b00001100, 8'b00000000, 8'b00000001, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10011010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 240: 
        // x=-98, 
        // s=[-1.  1. -1. -1.  1. -1. -1.  1.],
        // w=[ 6  0 10  2  0  5  1  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 10193. -12002.  34553.  22536. -27936. -19041.  49253. -40520.], 
        // Q{mac}=[ 9  0 33 22  0  0 48  0]

        sign=8'b01001001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000110, 8'b00000000, 8'b00001010, 8'b00000010, 8'b00000000, 8'b00000101, 8'b00000001, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10011110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 241: 
        // x=-101, 
        // s=[-1. -1.  1. -1.  1. -1.  1.  1.],
        // w=[ 6  6  4  5 13  6  6  8],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 10799. -11396.  34149.  23041. -29249. -18435.  48647. -41328.], 
        // Q{mac}=[10  0 33 22  0  0 47  0]

        sign=8'b00101011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000110, 8'b00000110, 8'b00000100, 8'b00000101, 8'b00001101, 8'b00000110, 8'b00000110, 8'b00001000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10011011;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 242: 
        // x=-92, 
        // s=[-1.  1. -1. -1. -1.  1. -1. -1.],
        // w=[ 1  3 14 14  3  1  1  1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 10891. -11672.  35437.  24329. -28973. -18527.  48739. -41236.], 
        // Q{mac}=[10  0 34 23  0  0 47  0]

        sign=8'b01000100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00000011, 8'b00001110, 8'b00001110, 8'b00000011, 8'b00000001, 8'b00000001, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10100100;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 243: 
        // x=-98, 
        // s=[-1.  1. -1. -1. -1.  1. -1.  1.],
        // w=[ 3  4  6 14  8 20  6 10],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 11185. -12064.  36025.  25701. -28189. -20487.  49327. -42216.], 
        // Q{mac}=[10  0 35 25  0  0 48  0]

        sign=8'b01000101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00000100, 8'b00000110, 8'b00001110, 8'b00001000, 8'b00010100, 8'b00000110, 8'b00001010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10011110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 244: 
        // x=-102, 
        // s=[-1. -1. -1. -1.  1.  1.  1. -1.],
        // w=[ 7  2  8 15  5  9  8  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 11899. -11860.  36841.  27231. -28699. -21405.  48511. -42012.], 
        // Q{mac}=[11  0 35 26  0  0 47  0]

        sign=8'b00001110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00000010, 8'b00001000, 8'b00001111, 8'b00000101, 8'b00001001, 8'b00001000, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10011010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 245: 
        // x=-125, 
        // s=[ 1. -1.  1. -1.  1. -1.  1.  1.],
        // w=[ 7  7  5 13  2  1  6  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 11024. -10985.  36216.  28856. -28949. -21280.  47761. -42387.], 
        // Q{mac}=[10  0 35 28  0  0 46  0]

        sign=8'b10101011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00000111, 8'b00000101, 8'b00001101, 8'b00000010, 8'b00000001, 8'b00000110, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000011;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 246: 
        // x=-108, 
        // s=[-1.  1.  1. -1.  1. -1. -1.  1.],
        // w=[2 7 8 1 8 5 1 5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 11240. -11741.  35352.  28964. -29813. -20740.  47869. -42927.], 
        // Q{mac}=[10  0 34 28  0  0 46  0]

        sign=8'b01101001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00000111, 8'b00001000, 8'b00000001, 8'b00001000, 8'b00000101, 8'b00000001, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10010100;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 247: 
        // x=84, 
        // s=[ 1.  1. -1.  1.  1.  1. -1.  1.],
        // w=[ 0  4 11  4  4 22  5  4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 11240. -11405.  34428.  29300. -29477. -18892.  47449. -42591.], 
        // Q{mac}=[10  0 33 28  0  0 46  0]

        sign=8'b11011101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000000, 8'b00000100, 8'b00001011, 8'b00000100, 8'b00000100, 8'b00010110, 8'b00000101, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b01010100;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 248: 
        // x=4, 
        // s=[ 1.  1. -1. -1.  1. -1. -1.  1.],
        // w=[ 3 16 16  1  8 12  5  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 11252. -11341.  34364.  29296. -29445. -18940.  47429. -42579.], 
        // Q{mac}=[10  0 33 28  0  0 46  0]

        sign=8'b11001001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00010000, 8'b00010000, 8'b00000001, 8'b00001000, 8'b00001100, 8'b00000101, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00000100;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 249: 
        // x=-22, 
        // s=[ 1. -1. -1. -1. -1.  1. -1. -1.],
        // w=[ 8  5  1 10  6 23  8  1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 11076. -11231.  34386.  29516. -29313. -19446.  47605. -42557.], 
        // Q{mac}=[10  0 33 28  0  0 46  0]

        sign=8'b10000100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001000, 8'b00000101, 8'b00000001, 8'b00001010, 8'b00000110, 8'b00010111, 8'b00001000, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11101010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 250: 
        // x=19, 
        // s=[-1.  1.  1.  1. -1. -1.  1.  1.],
        // w=[14  1 10  9  3  8 16  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 10810. -11212.  34576.  29687. -29370. -19598.  47909. -42500.], 
        // Q{mac}=[10  0 33 28  0  0 46  0]

        sign=8'b01110011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001110, 8'b00000001, 8'b00001010, 8'b00001001, 8'b00000011, 8'b00001000, 8'b00010000, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00010011;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 251: 
        // x=-2, 
        // s=[ 1. -1.  1.  1. -1.  1. -1.  1.],
        // w=[ 1 13 31  5  2 12 10  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 10808. -11186.  34514.  29677. -29366. -19622.  47929. -42504.], 
        // Q{mac}=[10  0 33 28  0  0 46  0]

        sign=8'b10110101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00001101, 8'b00011111, 8'b00000101, 8'b00000010, 8'b00001100, 8'b00001010, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11111110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 252: 
        // x=-119, 
        // s=[-1. -1.  1. -1. -1. -1. -1.  1.],
        // w=[3 8 5 4 4 2 7 1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 11165. -10234.  33919.  30153. -28890. -19384.  48762. -42623.], 
        // Q{mac}=[10  0 33 29  0  0 47  0]

        sign=8'b00100001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00001000, 8'b00000101, 8'b00000100, 8'b00000100, 8'b00000010, 8'b00000111, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 253: 
        // x=-115, 
        // s=[ 1.  1.  1.  1.  1. -1. -1.  1.],
        // w=[4 3 0 5 9 9 3 3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 10705. -10579.  33919.  29578. -29925. -18349.  49107. -42968.], 
        // Q{mac}=[10  0 33 28  0  0 47  0]

        sign=8'b11111001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000100, 8'b00000011, 8'b00000000, 8'b00000101, 8'b00001001, 8'b00001001, 8'b00000011, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 254: 
        // x=-116, 
        // s=[-1. -1. -1.  1. -1. -1. -1. -1.],
        // w=[7 5 4 2 4 2 4 2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 11517.  -9999.  34383.  29346. -29461. -18117.  49571. -42736.], 
        // Q{mac}=[11  0 33 28  0  0 48  0]

        sign=8'b00010000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00000101, 8'b00000100, 8'b00000010, 8'b00000100, 8'b00000010, 8'b00000100, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001100;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 255: 
        // x=-118, 
        // s=[-1. -1. -1. -1. -1.  1. -1. -1.],
        // w=[ 7  1  4 11  6  2  6  1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 12343.  -9881.  34855.  30644. -28753. -18353.  50279. -42618.], 
        // Q{mac}=[12  0 34 29  0  0 49  0]

        sign=8'b00000100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00000001, 8'b00000100, 8'b00001011, 8'b00000110, 8'b00000010, 8'b00000110, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 256: 
        // x=-125, 
        // s=[-1. -1.  1. -1. -1. -1. -1.  1.],
        // w=[15  6  8 10  4  3  1  6],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 14218.  -9131.  33855.  31894. -28253. -17978.  50404. -43368.], 
        // Q{mac}=[13  0 33 31  0  0 49  0]

        sign=8'b00100001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001111, 8'b00000110, 8'b00001000, 8'b00001010, 8'b00000100, 8'b00000011, 8'b00000001, 8'b00000110};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000011;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 257: 
        // x=-119, 
        // s=[-1. -1.  1. -1. -1. -1. -1.  1.],
        // w=[5 3 5 4 5 2 1 3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 14813.  -8774.  33260.  32370. -27658. -17740.  50523. -43725.], 
        // Q{mac}=[14  0 32 31  0  0 49  0]

        sign=8'b00100001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000101, 8'b00000011, 8'b00000101, 8'b00000100, 8'b00000101, 8'b00000010, 8'b00000001, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 258: 
        // x=-128, 
        // s=[-1.  1. -1.  1. -1.  1. -1.  1.],
        // w=[2 1 6 1 9 3 7 1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 15069.  -8902.  34028.  32242. -26506. -18124.  51419. -43853.], 
        // Q{mac}=[14  0 33 31  0  0 50  0]

        sign=8'b01010101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00000001, 8'b00000110, 8'b00000001, 8'b00001001, 8'b00000011, 8'b00000111, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 259: 
        // x=-117, 
        // s=[-1. -1.  1.  1.  1.  1. -1.  1.],
        // w=[11 11  9  5  2  5  8 10],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 16356.  -7615.  32975.  31657. -26740. -18709.  52355. -45023.], 
        // Q{mac}=[15  0 32 30  0  0 51  0]

        sign=8'b00111101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001011, 8'b00001011, 8'b00001001, 8'b00000101, 8'b00000010, 8'b00000101, 8'b00001000, 8'b00001010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001011;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 260: 
        // x=41, 
        // s=[-1.  1.  1. -1.  1. -1.  1. -1.],
        // w=[13  1  1  5 12  5  5  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 15823.  -7574.  33016.  31452. -26248. -18914.  52560. -45228.], 
        // Q{mac}=[15  0 32 30  0  0 51  0]

        sign=8'b01101010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001101, 8'b00000001, 8'b00000001, 8'b00000101, 8'b00001100, 8'b00000101, 8'b00000101, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00101001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 261: 
        // x=65, 
        // s=[ 1.  1.  1. -1. -1.  1.  1.  1.],
        // w=[ 0  9  4  3 20 23  4  0],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 15823.  -6989.  33276.  31257. -27548. -17419.  52820. -45228.], 
        // Q{mac}=[15  0 32 30  0  0 51  0]

        sign=8'b11100111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000000, 8'b00001001, 8'b00000100, 8'b00000011, 8'b00010100, 8'b00010111, 8'b00000100, 8'b00000000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b01000001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 262: 
        // x=-66, 
        // s=[-1.  1.  1. -1.  1. -1.  1. -1.],
        // w=[ 3  5  1  5 12 13  1  7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 16021.  -7319.  33210.  31587. -28340. -16561.  52754. -44766.], 
        // Q{mac}=[15  0 32 30  0  0 51  0]

        sign=8'b01101010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00000101, 8'b00000001, 8'b00000101, 8'b00001100, 8'b00001101, 8'b00000001, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10111110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 263: 
        // x=4, 
        // s=[-1. -1.  1. -1.  1. -1.  1. -1.],
        // w=[ 7 14  2  1 14 26  8  6],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 15993.  -7375.  33218.  31583. -28284. -16665.  52786. -44790.], 
        // Q{mac}=[15  0 32 30  0  0 51  0]

        sign=8'b00101010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00001110, 8'b00000010, 8'b00000001, 8'b00001110, 8'b00011010, 8'b00001000, 8'b00000110};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00000100;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 264: 
        // x=1, 
        // s=[ 1.  1.  1.  1. -1.  1. -1. -1.],
        // w=[18 11  3 12 14  4 22  9],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 16011.  -7364.  33221.  31595. -28298. -16661.  52764. -44799.], 
        // Q{mac}=[15  0 32 30  0  0 51  0]

        sign=8'b11110100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00010010, 8'b00001011, 8'b00000011, 8'b00001100, 8'b00001110, 8'b00000100, 8'b00010110, 8'b00001001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00000001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 265: 
        // x=-118, 
        // s=[-1.  1. -1. -1. -1.  1.  1. -1.],
        // w=[ 7 14 12 19  8 13  9  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 16837.  -9016.  34637.  33837. -27354. -18195.  51702. -44563.], 
        // Q{mac}=[16  0 33 33  0  0 50  0]

        sign=8'b01000110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00001110, 8'b00001100, 8'b00010011, 8'b00001000, 8'b00001101, 8'b00001001, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 266: 
        // x=-118, 
        // s=[-1. -1.  1. -1.  1.  1.  1.  1.],
        // w=[ 4 11  2  6 10  8  2  9],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 17309.  -7718.  34401.  34545. -28534. -19139.  51466. -45625.], 
        // Q{mac}=[16  0 33 33  0  0 50  0]

        sign=8'b00101111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000100, 8'b00001011, 8'b00000010, 8'b00000110, 8'b00001010, 8'b00001000, 8'b00000010, 8'b00001001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 267: 
        // x=-102, 
        // s=[-1. -1. -1. -1.  1.  1. -1.  1.],
        // w=[ 1  5  7 10  2  3  6  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 17411.  -7208.  35115.  35565. -28738. -19445.  52078. -45829.], 
        // Q{mac}=[17  0 34 34  0  0 50  0]

        sign=8'b00001101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00000101, 8'b00000111, 8'b00001010, 8'b00000010, 8'b00000011, 8'b00000110, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10011010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 268: 
        // x=-122, 
        // s=[ 1.  1. -1. -1. -1.  1.  1. -1.],
        // w=[ 1  5 14 26  6 15 13  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 17289.  -7818.  36823.  38737. -28006. -21275.  50492. -45463.], 
        // Q{mac}=[16  0 35 37  0  0 49  0]

        sign=8'b11000110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00000101, 8'b00001110, 8'b00011010, 8'b00000110, 8'b00001111, 8'b00001101, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 269: 
        // x=-119, 
        // s=[-1. -1.  1. -1.  1.  1.  1.  1.],
        // w=[ 9 13  6  3  2 18  3  0],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 18360.  -6271.  36109.  39094. -28244. -23417.  50135. -45463.], 
        // Q{mac}=[17  0 35 38  0  0 48  0]

        sign=8'b00101111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001001, 8'b00001101, 8'b00000110, 8'b00000011, 8'b00000010, 8'b00010010, 8'b00000011, 8'b00000000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 270: 
        // x=-82, 
        // s=[-1. -1.  1. -1.  1.  1.  1. -1.],
        // w=[ 5  7 11  3  0  6  3  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 18770.  -5697.  35207.  39340. -28244. -23909.  49889. -45299.], 
        // Q{mac}=[18  0 34 38  0  0 48  0]

        sign=8'b00101110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000101, 8'b00000111, 8'b00001011, 8'b00000011, 8'b00000000, 8'b00000110, 8'b00000011, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10101110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 271: 
        // x=-120, 
        // s=[-1.  1. -1. -1. -1.  1.  1.  1.],
        // w=[ 5  6 11 21  5 16  6  8],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 19370.  -6417.  36527.  41860. -27644. -25829.  49169. -46259.], 
        // Q{mac}=[18  0 35 40  0  0 48  0]

        sign=8'b01000111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000101, 8'b00000110, 8'b00001011, 8'b00010101, 8'b00000101, 8'b00010000, 8'b00000110, 8'b00001000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 272: 
        // x=-119, 
        // s=[-1. -1. -1.  1.  1.  1.  1.  1.],
        // w=[ 9  9  2  4  8 13  3 10],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 20441.  -5346.  36765.  41384. -28596. -27376.  48812. -47449.], 
        // Q{mac}=[19  0 35 40  0  0 47  0]

        sign=8'b00011111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001001, 8'b00001001, 8'b00000010, 8'b00000100, 8'b00001000, 8'b00001101, 8'b00000011, 8'b00001010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 273: 
        // x=-93, 
        // s=[-1.  1. -1. -1.  1.  1. -1. -1.],
        // w=[16  4  1  2  8  0  2  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 21929.  -5718.  36858.  41570. -29340. -27376.  48998. -47170.], 
        // Q{mac}=[21  0 35 40  0  0 47  0]

        sign=8'b01001100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00010000, 8'b00000100, 8'b00000001, 8'b00000010, 8'b00001000, 8'b00000000, 8'b00000010, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10100011;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 274: 
        // x=-124, 
        // s=[ 1.  1. -1. -1. -1.  1.  1.  1.],
        // w=[14 13 12 26  2 18  9 10],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 20193.  -7330.  38346.  44794. -29092. -29608.  47882. -48410.], 
        // Q{mac}=[19  0 37 43  0  0 46  0]

        sign=8'b11000111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001110, 8'b00001101, 8'b00001100, 8'b00011010, 8'b00000010, 8'b00010010, 8'b00001001, 8'b00001010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000100;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 275: 
        // x=-121, 
        // s=[-1. -1.  1.  1. -1.  1.  1.  1.],
        // w=[ 6  4  4  8 14 10  6  0],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 20919.  -6846.  37862.  43826. -27398. -30818.  47156. -48410.], 
        // Q{mac}=[20  0 36 42  0  0 46  0]

        sign=8'b00110111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000110, 8'b00000100, 8'b00000100, 8'b00001000, 8'b00001110, 8'b00001010, 8'b00000110, 8'b00000000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000111;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 276: 
        // x=-77, 
        // s=[ 1. -1.  1.  1. -1. -1. -1. -1.],
        // w=[ 2  7  9  1 11  2  4  6],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 20765.  -6307.  37169.  43749. -26551. -30664.  47464. -47948.], 
        // Q{mac}=[20  0 36 42  0  0 46  0]

        sign=8'b10110000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00000111, 8'b00001001, 8'b00000001, 8'b00001011, 8'b00000010, 8'b00000100, 8'b00000110};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10110011;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 277: 
        // x=-124, 
        // s=[ 1. -1. -1.  1. -1.  1. -1.  1.],
        // w=[1 2 3 1 1 5 7 1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 20641.  -6059.  37541.  43625. -26427. -31284.  48332. -48072.], 
        // Q{mac}=[20  0 36 42  0  0 47  0]

        sign=8'b10010101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00000010, 8'b00000011, 8'b00000001, 8'b00000001, 8'b00000101, 8'b00000111, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000100;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 278: 
        // x=-127, 
        // s=[ 1. -1. -1. -1.  1.  1. -1.  1.],
        // w=[7 6 6 2 3 0 8 5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 19752.  -5297.  38303.  43879. -26808. -31284.  49348. -48707.], 
        // Q{mac}=[19  0 37 42  0  0 48  0]

        sign=8'b10001101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00000110, 8'b00000110, 8'b00000010, 8'b00000011, 8'b00000000, 8'b00001000, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 279: 
        // x=-122, 
        // s=[-1. -1. -1.  1.  1.  1. -1.  1.],
        // w=[3 2 6 1 1 1 4 9],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 20118.  -5053.  39035.  43757. -26930. -31406.  49836. -49805.], 
        // Q{mac}=[19  0 38 42  0  0 48  0]

        sign=8'b00011101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00000010, 8'b00000110, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000100, 8'b00001001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 280: 
        // x=-111, 
        // s=[-1.  1. -1. -1.  1.  1. -1.  1.],
        // w=[ 1 12  9  1 13 11  1  6],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 20229.  -6385.  40034.  43868. -28373. -32627.  49947. -50471.], 
        // Q{mac}=[19  0 39 42  0  0 48  0]

        sign=8'b01001101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00001100, 8'b00001001, 8'b00000001, 8'b00001101, 8'b00001011, 8'b00000001, 8'b00000110};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10010001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 281: 
        // x=-128, 
        // s=[ 1.  1. -1. -1. -1.  1.  1.  1.],
        // w=[ 4  1  6 10  2  8  6  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 19717.  -6513.  40802.  45148. -28117. -33651.  49179. -51111.], 
        // Q{mac}=[19  0 39 44  0  0 48  0]

        sign=8'b11000111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000100, 8'b00000001, 8'b00000110, 8'b00001010, 8'b00000010, 8'b00001000, 8'b00000110, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 282: 
        // x=-128, 
        // s=[-1. -1.  1.  1. -1.  1.  1.  1.],
        // w=[ 1 11  5  0  6  8  4  7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 19845.  -5105.  40162.  45148. -27349. -34675.  48667. -52007.], 
        // Q{mac}=[19  0 39 44  0  0 47  0]

        sign=8'b00110111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00001011, 8'b00000101, 8'b00000000, 8'b00000110, 8'b00001000, 8'b00000100, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 283: 
        // x=-121, 
        // s=[ 1. -1. -1. -1.  1. -1. -1. -1.],
        // w=[0 4 2 4 1 6 1 4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 19845.  -4621.  40404.  45632. -27470. -33949.  48788. -51523.], 
        // Q{mac}=[19  0 39 44  0  0 47  0]

        sign=8'b10001000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000000, 8'b00000100, 8'b00000010, 8'b00000100, 8'b00000001, 8'b00000110, 8'b00000001, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000111;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 284: 
        // x=-116, 
        // s=[-1.  1. -1. -1. -1.  1.  1.  1.],
        // w=[13 10  4 16  2  8 10  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 21353.  -5781.  40868.  47488. -27238. -34877.  47628. -52103.], 
        // Q{mac}=[20  0 39 46  0  0 46  0]

        sign=8'b01000111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001101, 8'b00001010, 8'b00000100, 8'b00010000, 8'b00000010, 8'b00001000, 8'b00001010, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001100;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 285: 
        // x=-120, 
        // s=[-1. -1.  1.  1.  1.  1.  1. -1.],
        // w=[2 8 0 0 2 0 9 2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 21593.  -4821.  40868.  47488. -27478. -34877.  46548. -51863.], 
        // Q{mac}=[21  0 39 46  0  0 45  0]

        sign=8'b00111110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00001000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000000, 8'b00001001, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 286: 
        // x=-112, 
        // s=[-1.  1. -1. -1.  1.  1.  1. -1.],
        // w=[10  2  1  9 18  1  5  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 22713.  -5045.  40980.  48496. -29494. -34989.  45988. -51639.], 
        // Q{mac}=[22  0 40 47  0  0 44  0]

        sign=8'b01001110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001010, 8'b00000010, 8'b00000001, 8'b00001001, 8'b00010010, 8'b00000001, 8'b00000101, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10010000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 287: 
        // x=-44, 
        // s=[-1.  1. -1. -1.  1.  1.  1. -1.],
        // w=[13  4 11 11  8  4  7  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 23285.  -5221.  41464.  48980. -29846. -35165.  45680. -51419.], 
        // Q{mac}=[22  0 40 47  0  0 44  0]

        sign=8'b01001110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001101, 8'b00000100, 8'b00001011, 8'b00001011, 8'b00001000, 8'b00000100, 8'b00000111, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11010100;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 288: 
        // x=-63, 
        // s=[-1.  1. -1. -1.  1.  1.  1.  1.],
        // w=[ 3  2  9  9 23 14  8  0],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 23474.  -5347.  42031.  49547. -31295. -36047.  45176. -51419.], 
        // Q{mac}=[22  0 41 48  0  0 44  0]

        sign=8'b01001111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00000010, 8'b00001001, 8'b00001001, 8'b00010111, 8'b00001110, 8'b00001000, 8'b00000000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11000001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 289: 
        // x=-22, 
        // s=[-1.  1. -1. -1.  1. -1.  1.  1.],
        // w=[ 7  6  9  4 31  1  2  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 23628.  -5479.  42229.  49635. -31977. -36025.  45132. -51529.], 
        // Q{mac}=[23  0 41 48  0  0 44  0]

        sign=8'b01001011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00000110, 8'b00001001, 8'b00000100, 8'b00011111, 8'b00000001, 8'b00000010, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11101010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 290: 
        // x=-128, 
        // s=[ 1. -1. -1.  1. -1.  1. -1. -1.],
        // w=[ 1  3  4  1  4  6 13  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 23500.  -5095.  42741.  49507. -31465. -36793.  46796. -51145.], 
        // Q{mac}=[22  0 41 48  0  0 45  0]

        sign=8'b10010100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00000011, 8'b00000100, 8'b00000001, 8'b00000100, 8'b00000110, 8'b00001101, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 291: 
        // x=-128, 
        // s=[ 1.  1. -1. -1.  1. -1. -1.  1.],
        // w=[ 7  7  3  4 11  7 16  6],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 22604.  -5991.  43125.  50019. -32873. -35897.  48844. -51913.], 
        // Q{mac}=[22  0 42 48  0  0 47  0]

        sign=8'b11001001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00000111, 8'b00000011, 8'b00000100, 8'b00001011, 8'b00000111, 8'b00010000, 8'b00000110};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 292: 
        // x=-128, 
        // s=[ 1.  1. -1. -1.  1. -1. -1.  1.],
        // w=[ 3  5  1  5  0  3 11  6],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 22220.  -6631.  43253.  50659. -32873. -35513.  50252. -52681.], 
        // Q{mac}=[21  0 42 49  0  0 49  0]

        sign=8'b11001001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00000101, 8'b00000001, 8'b00000101, 8'b00000000, 8'b00000011, 8'b00001011, 8'b00000110};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 293: 
        // x=14, 
        // s=[-1. -1. -1.  1.  1. -1. -1.  1.],
        // w=[ 7  3  4  0 38 25 13  7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 22122.  -6673.  43197.  50659. -32341. -35863.  50070. -52583.], 
        // Q{mac}=[21  0 42 49  0  0 48  0]

        sign=8'b00011001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00000011, 8'b00000100, 8'b00000000, 8'b00100110, 8'b00011001, 8'b00001101, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00001110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 294: 
        // x=-68, 
        // s=[-1. -1. -1.  1.  1. -1.  1.  1.],
        // w=[ 9  2 21 15 33 32 10  6],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 22734.  -6537.  44625.  49639. -34585. -33687.  49390. -52991.], 
        // Q{mac}=[22  0 43 48  0  0 48  0]

        sign=8'b00011011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001001, 8'b00000010, 8'b00010101, 8'b00001111, 8'b00100001, 8'b00100000, 8'b00001010, 8'b00000110};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10111100;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 295: 
        // x=-74, 
        // s=[ 1.  1. -1. -1. -1.  1. -1. -1.],
        // w=[21 10  1 30 11 27  3  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 21180.  -7277.  44699.  51859. -33771. -35685.  49612. -52843.], 
        // Q{mac}=[20  0 43 50  0  0 48  0]

        sign=8'b11000100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00010101, 8'b00001010, 8'b00000001, 8'b00011110, 8'b00001011, 8'b00011011, 8'b00000011, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10110110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 296: 
        // x=-115, 
        // s=[ 1.  1. -1. -1. -1.  1. -1.  1.],
        // w=[20  4  4 17 17 24  2 10],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 18880.  -7737.  45159.  53814. -31816. -38445.  49842. -53993.], 
        // Q{mac}=[18  0 44 52  0  0 48  0]

        sign=8'b11000101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00010100, 8'b00000100, 8'b00000100, 8'b00010001, 8'b00010001, 8'b00011000, 8'b00000010, 8'b00001010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 297: 
        // x=-44, 
        // s=[ 1. -1.  1.  1. -1.  1.  1.  1.],
        // w=[ 3 21  9 30 25  7 15  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 18748.  -6813.  44763.  52494. -30716. -38753.  49182. -54081.], 
        // Q{mac}=[18  0 43 51  0  0 48  0]

        sign=8'b10110111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00010101, 8'b00001001, 8'b00011110, 8'b00011001, 8'b00000111, 8'b00001111, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11010100;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 298: 
        // x=-89, 
        // s=[-1. -1.  1.  1. -1. -1.  1.  1.],
        // w=[ 1 21  0 18 21  3  1  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 18837.  -4944.  44763.  50892. -28847. -38486.  49093. -54348.], 
        // Q{mac}=[18  0 43 49  0  0 47  0]

        sign=8'b00110011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00010101, 8'b00000000, 8'b00010010, 8'b00010101, 8'b00000011, 8'b00000001, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10100111;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 299: 
        // x=23, 
        // s=[ 1. -1.  1.  1. -1. -1.  1.  1.],
        // w=[ 1 11  7 11  9 15  0  1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 18860.  -5197.  44924.  51145. -29054. -38831.  49093. -54325.], 
        // Q{mac}=[18  0 43 49  0  0 47  0]

        sign=8'b10110011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00001011, 8'b00000111, 8'b00001011, 8'b00001001, 8'b00001111, 8'b00000000, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00010111;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 300: 
        // x=-15, 
        // s=[ 1. -1.  1.  1. -1. -1.  1. -1.],
        // w=[10 16  0  5 14 12  5  1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 18710.  -4957.  44924.  51070. -28844. -38651.  49018. -54310.], 
        // Q{mac}=[18  0 43 49  0  0 47  0]

        sign=8'b10110010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001010, 8'b00010000, 8'b00000000, 8'b00000101, 8'b00001110, 8'b00001100, 8'b00000101, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11110001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 301: 
        // x=-128, 
        // s=[ 1.  1. -1. -1. -1.  1.  1.  1.],
        // w=[ 1  6  7 11  2 10  2  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 18582.  -5725.  45820.  52478. -28588. -39931.  48762. -54694.], 
        // Q{mac}=[18  0 44 51  0  0 47  0]

        sign=8'b11000111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00000110, 8'b00000111, 8'b00001011, 8'b00000010, 8'b00001010, 8'b00000010, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 302: 
        // x=-128, 
        // s=[-1.  1. -1. -1. -1.  1.  1.  1.],
        // w=[1 5 3 6 2 6 0 6],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 18710.  -6365.  46204.  53246. -28332. -40699.  48762. -55462.], 
        // Q{mac}=[18  0 45 51  0  0 47  0]

        sign=8'b01000111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00000101, 8'b00000011, 8'b00000110, 8'b00000010, 8'b00000110, 8'b00000000, 8'b00000110};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 303: 
        // x=-128, 
        // s=[-1.  1.  1. -1.  1. -1. -1.  1.],
        // w=[1 4 2 7 4 1 6 0],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 18838.  -6877.  45948.  54142. -28844. -40571.  49530. -55462.], 
        // Q{mac}=[18  0 44 52  0  0 48  0]

        sign=8'b01101001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00000100, 8'b00000010, 8'b00000111, 8'b00000100, 8'b00000001, 8'b00000110, 8'b00000000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 304: 
        // x=-128, 
        // s=[-1. -1. -1. -1.  1.  1.  1.  1.],
        // w=[1 4 4 8 0 3 3 3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 18966.  -6365.  46460.  55166. -28844. -40955.  49146. -55846.], 
        // Q{mac}=[18  0 45 53  0  0 47  0]

        sign=8'b00001111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00000100, 8'b00000100, 8'b00001000, 8'b00000000, 8'b00000011, 8'b00000011, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 305: 
        // x=-128, 
        // s=[-1.  1. -1. -1. -1. -1. -1.  1.],
        // w=[5 1 3 2 3 4 7 6],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 19606.  -6493.  46844.  55422. -28460. -40443.  50042. -56614.], 
        // Q{mac}=[19  0 45 54  0  0 48  0]

        sign=8'b01000001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000101, 8'b00000001, 8'b00000011, 8'b00000010, 8'b00000011, 8'b00000100, 8'b00000111, 8'b00000110};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 306: 
        // x=-127, 
        // s=[ 1.  1.  1. -1. -1.  1.  1.  1.],
        // w=[ 0 11  2  5  8  9  1  1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 19606.  -7890.  46590.  56057. -27444. -41586.  49915. -56741.], 
        // Q{mac}=[19  0 45 54  0  0 48  0]

        sign=8'b11100111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000000, 8'b00001011, 8'b00000010, 8'b00000101, 8'b00001000, 8'b00001001, 8'b00000001, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 307: 
        // x=-127, 
        // s=[-1. -1.  1. -1.  1. -1. -1.  1.],
        // w=[4 4 3 8 2 7 7 1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 20114.  -7382.  46209.  57073. -27698. -40697.  50804. -56868.], 
        // Q{mac}=[19  0 45 55  0  0 49  0]

        sign=8'b00101001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000100, 8'b00000100, 8'b00000011, 8'b00001000, 8'b00000010, 8'b00000111, 8'b00000111, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 308: 
        // x=-128, 
        // s=[ 1. -1.  1. -1.  1.  1.  1. -1.],
        // w=[5 1 1 2 1 4 3 1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 19474.  -7254.  46081.  57329. -27826. -41209.  50420. -56740.], 
        // Q{mac}=[19  0 45 55  0  0 49  0]

        sign=8'b10101110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000101, 8'b00000001, 8'b00000001, 8'b00000010, 8'b00000001, 8'b00000100, 8'b00000011, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 309: 
        // x=-128, 
        // s=[ 1.  1. -1. -1. -1.  1. -1.  1.],
        // w=[ 2 16  8 10  5 10  3  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 19218.  -9302.  47105.  58609. -27186. -42489.  50804. -57380.], 
        // Q{mac}=[18  0 46 57  0  0 49  0]

        sign=8'b11000101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00010000, 8'b00001000, 8'b00001010, 8'b00000101, 8'b00001010, 8'b00000011, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 310: 
        // x=-128, 
        // s=[-1. -1.  1. -1. -1. -1. -1. -1.],
        // w=[7 5 0 4 9 5 6 1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 20114.  -8662.  47105.  59121. -26034. -41849.  51572. -57252.], 
        // Q{mac}=[19  0 46 57  0  0 50  0]

        sign=8'b00100000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00000101, 8'b00000000, 8'b00000100, 8'b00001001, 8'b00000101, 8'b00000110, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 311: 
        // x=-128, 
        // s=[-1. -1. -1. -1. -1. -1.  1.  1.],
        // w=[2 4 3 8 9 1 6 2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 20370.  -8150.  47489.  60145. -24882. -41721.  50804. -57508.], 
        // Q{mac}=[19  0 46 58  0  0 49  0]

        sign=8'b00000011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00000100, 8'b00000011, 8'b00001000, 8'b00001001, 8'b00000001, 8'b00000110, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 312: 
        // x=-128, 
        // s=[ 1. -1. -1. -1. -1. -1.  1. -1.],
        // w=[8 4 7 5 3 3 7 1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 19346.  -7638.  48385.  60785. -24498. -41337.  49908. -57380.], 
        // Q{mac}=[18  0 47 59  0  0 48  0]

        sign=8'b10000010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001000, 8'b00000100, 8'b00000111, 8'b00000101, 8'b00000011, 8'b00000011, 8'b00000111, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 313: 
        // x=-128, 
        // s=[ 1.  1. -1. -1.  1.  1.  1.  1.],
        // w=[11 14 14  4  4  5  5  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 17938.  -9430.  50177.  61297. -25010. -41977.  49268. -57764.], 
        // Q{mac}=[17  0 49 59  0  0 48  0]

        sign=8'b11001111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001011, 8'b00001110, 8'b00001110, 8'b00000100, 8'b00000100, 8'b00000101, 8'b00000101, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 314: 
        // x=-128, 
        // s=[-1.  1. -1. -1. -1. -1.  1.  1.],
        // w=[ 4  3 10  8  8  4  0  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 18450.  -9814.  51457.  62321. -23986. -41465.  49268. -58404.], 
        // Q{mac}=[18  0 50 60  0  0 48  0]

        sign=8'b01000011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000100, 8'b00000011, 8'b00001010, 8'b00001000, 8'b00001000, 8'b00000100, 8'b00000000, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 315: 
        // x=-128, 
        // s=[-1. -1.  1.  1. -1.  1.  1.  1.],
        // w=[ 1  1  1  6 12 17  2  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 18578.  -9686.  51329.  61553. -22450. -43641.  49012. -59044.], 
        // Q{mac}=[18  0 50 60  0  0 47  0]

        sign=8'b00110111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00000001, 8'b00000001, 8'b00000110, 8'b00001100, 8'b00010001, 8'b00000010, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 316: 
        // x=-128, 
        // s=[-1. -1.  1.  1. -1. -1.  1.  1.],
        // w=[4 4 6 9 1 3 2 2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 19090.  -9174.  50561.  60401. -22322. -43257.  48756. -59300.], 
        // Q{mac}=[18  0 49 58  0  0 47  0]

        sign=8'b00110011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000100, 8'b00000100, 8'b00000110, 8'b00001001, 8'b00000001, 8'b00000011, 8'b00000010, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 317: 
        // x=-128, 
        // s=[-1. -1.  1.  1. -1. -1.  1.  1.],
        // w=[9 5 6 2 4 1 7 7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 20242.  -8534.  49793.  60145. -21810. -43129.  47860. -60196.], 
        // Q{mac}=[19  0 48 58  0  0 46  0]

        sign=8'b00110011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001001, 8'b00000101, 8'b00000110, 8'b00000010, 8'b00000100, 8'b00000001, 8'b00000111, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 318: 
        // x=-128, 
        // s=[ 1.  1. -1. -1. -1. -1. -1. -1.],
        // w=[3 4 1 5 5 7 3 2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 19858.  -9046.  49921.  60785. -21170. -42233.  48244. -59940.], 
        // Q{mac}=[19  0 48 59  0  0 47  0]

        sign=8'b11000000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00000100, 8'b00000001, 8'b00000101, 8'b00000101, 8'b00000111, 8'b00000011, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 319: 
        // x=-128, 
        // s=[ 1. -1. -1.  1. -1. -1. -1.  1.],
        // w=[3 1 3 0 5 8 3 4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 19474.  -8918.  50305.  60785. -20530. -41209.  48628. -60452.], 
        // Q{mac}=[19  0 49 59  0  0 47  0]

        sign=8'b10010001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00000001, 8'b00000011, 8'b00000000, 8'b00000101, 8'b00001000, 8'b00000011, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 320: 
        // x=-128, 
        // s=[-1. -1.  1. -1. -1. -1. -1. -1.],
        // w=[8 3 2 7 9 4 8 4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 20498.  -8534.  50049.  61681. -19378. -40697.  49652. -59940.], 
        // Q{mac}=[20  0 48 60  0  0 48  0]

        sign=8'b00100000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001000, 8'b00000011, 8'b00000010, 8'b00000111, 8'b00001001, 8'b00000100, 8'b00001000, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 321: 
        // x=-128, 
        // s=[-1. -1. -1. -1. -1. -1. -1. -1.],
        // w=[ 2  8  1  7  3 10  6  1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 20754.  -7510.  50177.  62577. -18994. -39417.  50420. -59812.], 
        // Q{mac}=[20  0 49 61  0  0 49  0]

        sign=8'b00000000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00001000, 8'b00000001, 8'b00000111, 8'b00000011, 8'b00001010, 8'b00000110, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 322: 
        // x=-128, 
        // s=[ 1.  1. -1. -1.  1. -1. -1. -1.],
        // w=[7 2 8 6 4 3 2 3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 19858.  -7766.  51201.  63345. -19506. -39033.  50676. -59428.], 
        // Q{mac}=[19  0 50 61  0  0 49  0]

        sign=8'b11001000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00000010, 8'b00001000, 8'b00000110, 8'b00000100, 8'b00000011, 8'b00000010, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 323: 
        // x=-128, 
        // s=[-1. -1.  1.  1. -1.  1. -1.  1.],
        // w=[7 2 1 0 2 1 2 7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 20754.  -7510.  51073.  63345. -19250. -39161.  50932. -60324.], 
        // Q{mac}=[20  0 49 61  0  0 49  0]

        sign=8'b00110101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000010, 8'b00000001, 8'b00000010, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 324: 
        // x=-128, 
        // s=[-1. -1.  1.  1. -1.  1. -1.  1.],
        // w=[ 3  9  7  7 10  3  6  7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 21138.  -6358.  50177.  62449. -17970. -39545.  51700. -61220.], 
        // Q{mac}=[20  0 49 60  0  0 50  0]

        sign=8'b00110101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00001001, 8'b00000111, 8'b00000111, 8'b00001010, 8'b00000011, 8'b00000110, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 325: 
        // x=-128, 
        // s=[ 1. -1.  1. -1.  1. -1. -1. -1.],
        // w=[3 5 2 5 1 1 7 4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 20754.  -5718.  49921.  63089. -18098. -39417.  52596. -60708.], 
        // Q{mac}=[20  0 48 61  0  0 51  0]

        sign=8'b10101000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00000101, 8'b00000010, 8'b00000101, 8'b00000001, 8'b00000001, 8'b00000111, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 326: 
        // x=-128, 
        // s=[ 1.  1. -1. -1. -1. -1. -1. -1.],
        // w=[3 6 4 2 6 2 5 6],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 20370.  -6486.  50433.  63345. -17330. -39161.  53236. -59940.], 
        // Q{mac}=[19  0 49 61  0  0 51  0]

        sign=8'b11000000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00000110, 8'b00000100, 8'b00000010, 8'b00000110, 8'b00000010, 8'b00000101, 8'b00000110};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 327: 
        // x=-128, 
        // s=[-1. -1. -1.  1. -1.  1. -1.  1.],
        // w=[ 3 10  2  5  1  2  6  0],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 20754.  -5206.  50689.  62705. -17202. -39417.  54004. -59940.], 
        // Q{mac}=[20  0 49 61  0  0 52  0]

        sign=8'b00010101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00001010, 8'b00000010, 8'b00000101, 8'b00000001, 8'b00000010, 8'b00000110, 8'b00000000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 328: 
        // x=-128, 
        // s=[ 1. -1. -1.  1.  1.  1.  1.  1.],
        // w=[ 1 10  1  7  7  1  3  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 20626.  -3926.  50817.  61809. -18098. -39545.  53620. -60580.], 
        // Q{mac}=[20  0 49 60  0  0 52  0]

        sign=8'b10011111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00001010, 8'b00000001, 8'b00000111, 8'b00000111, 8'b00000001, 8'b00000011, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 329: 
        // x=-119, 
        // s=[-1. -1.  1. -1. -1. -1. -1.  1.],
        // w=[ 9 10  4  5  3  4  8  1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 21697.  -2736.  50341.  62404. -17741. -39069.  54572. -60699.], 
        // Q{mac}=[21  0 49 60  0  0 53  0]

        sign=8'b00100001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001001, 8'b00001010, 8'b00000100, 8'b00000101, 8'b00000011, 8'b00000100, 8'b00001000, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 330: 
        // x=-128, 
        // s=[ 1.  1.  1. -1. -1. -1. -1.  1.],
        // w=[2 4 5 7 4 7 7 3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 21441.  -3248.  49701.  63300. -17229. -38173.  55468. -61083.], 
        // Q{mac}=[20  0 48 61  0  0 54  0]

        sign=8'b11100001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00000100, 8'b00000101, 8'b00000111, 8'b00000100, 8'b00000111, 8'b00000111, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 331: 
        // x=-128, 
        // s=[ 1.  1. -1.  1.  1. -1. -1.  1.],
        // w=[ 1  1  9  0  2  4 10  4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 21313.  -3376.  50853.  63300. -17485. -37661.  56748. -61595.], 
        // Q{mac}=[20  0 49 61  0  0 55  0]

        sign=8'b11011001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00000001, 8'b00001001, 8'b00000000, 8'b00000010, 8'b00000100, 8'b00001010, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 332: 
        // x=-128, 
        // s=[ 1. -1.  1. -1. -1.  1. -1.  1.],
        // w=[6 1 3 7 6 1 2 7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 20545.  -3248.  50469.  64196. -16717. -37789.  57004. -62491.], 
        // Q{mac}=[20  0 49 62  0  0 55  0]

        sign=8'b10100101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000110, 8'b00000001, 8'b00000011, 8'b00000111, 8'b00000110, 8'b00000001, 8'b00000010, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 333: 
        // x=-128, 
        // s=[-1.  1.  1. -1. -1.  1. -1.  1.],
        // w=[5 1 0 9 4 1 4 7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 21185.  -3376.  50469.  65348. -16205. -37917.  57516. -63387.], 
        // Q{mac}=[20  0 49 63  0  0 56  0]

        sign=8'b01100101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000101, 8'b00000001, 8'b00000000, 8'b00001001, 8'b00000100, 8'b00000001, 8'b00000100, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 334: 
        // x=-128, 
        // s=[-1.  1. -1.  1. -1. -1.  1.  1.],
        // w=[9 3 5 2 6 5 4 8],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 22337.  -3760.  51109.  65092. -15437. -37277.  57004. -64411.], 
        // Q{mac}=[21  0 49 63  0  0 55  0]

        sign=8'b01010011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001001, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000110, 8'b00000101, 8'b00000100, 8'b00001000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 335: 
        // x=-127, 
        // s=[ 1.  1. -1.  1. -1. -1.  1. -1.],
        // w=[0 2 4 0 4 6 5 1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 22337.  -4014.  51617.  65092. -14929. -36515.  56369. -64284.], 
        // Q{mac}=[21  0 50 63  0  0 55  0]

        sign=8'b11010010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000000, 8'b00000010, 8'b00000100, 8'b00000000, 8'b00000100, 8'b00000110, 8'b00000101, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 336: 
        // x=-126, 
        // s=[-1. -1.  1.  1. -1.  1. -1. -1.],
        // w=[ 2  4  3  0 12  7  9  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 22589.  -3510.  51239.  65092. -13417. -37397.  57503. -64032.], 
        // Q{mac}=[22  0 50 63  0  0 56  0]

        sign=8'b00110100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00000100, 8'b00000011, 8'b00000000, 8'b00001100, 8'b00000111, 8'b00001001, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 337: 
        // x=-121, 
        // s=[-1.  1.  1. -1. -1. -1. -1. -1.],
        // w=[8 2 3 2 5 1 5 3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 23557.  -3752.  50876.  65334. -12812. -37276.  58108. -63669.], 
        // Q{mac}=[23  0 49 63  0  0 56  0]

        sign=8'b01100000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001000, 8'b00000010, 8'b00000011, 8'b00000010, 8'b00000101, 8'b00000001, 8'b00000101, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000111;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 338: 
        // x=-128, 
        // s=[-1.  1. -1.  1.  1. -1. -1. -1.],
        // w=[8 7 4 4 9 6 5 1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 24581.  -4648.  51388.  64822. -13964. -36508.  58748. -63541.], 
        // Q{mac}=[24  0 50 63  0  0 57  0]

        sign=8'b01011000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001000, 8'b00000111, 8'b00000100, 8'b00000100, 8'b00001001, 8'b00000110, 8'b00000101, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 339: 
        // x=-128, 
        // s=[-1. -1. -1.  1. -1. -1. -1. -1.],
        // w=[ 8  8  3  2  4 10 10  4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 25605.  -3624.  51772.  64566. -13452. -35228.  60028. -63029.], 
        // Q{mac}=[25  0 50 63  0  0 58  0]

        sign=8'b00010000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001000, 8'b00001000, 8'b00000011, 8'b00000010, 8'b00000100, 8'b00001010, 8'b00001010, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 340: 
        // x=-127, 
        // s=[-1. -1. -1. -1.  1.  1.  1.  1.],
        // w=[2 8 8 9 0 1 4 9],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 25859.  -2608.  52788.  65709. -13452. -35355.  59520. -64172.], 
        // Q{mac}=[25  0 51 64  0  0 58  0]

        sign=8'b00001111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00001000, 8'b00001000, 8'b00001001, 8'b00000000, 8'b00000001, 8'b00000100, 8'b00001001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 341: 
        // x=-121, 
        // s=[ 1.  1. -1.  1. -1. -1.  1.  1.],
        // w=[2 4 6 6 4 4 6 2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 25617.  -3092.  53514.  64983. -12968. -34871.  58794. -64414.], 
        // Q{mac}=[25  0 52 63  0  0 57  0]

        sign=8'b11010011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00000100, 8'b00000110, 8'b00000110, 8'b00000100, 8'b00000100, 8'b00000110, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000111;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 342: 
        // x=-128, 
        // s=[-1. -1.  1. -1. -1.  1.  1.  1.],
        // w=[7 7 0 7 2 2 1 8],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 26513.  -2196.  53514.  65879. -12712. -35127.  58666. -65438.], 
        // Q{mac}=[25  0 52 64  0  0 57  0]

        sign=8'b00100111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00000111, 8'b00000000, 8'b00000111, 8'b00000010, 8'b00000010, 8'b00000001, 8'b00001000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 343: 
        // x=-116, 
        // s=[-1.  1. -1. -1.  1.  1.  1.  1.],
        // w=[ 9  8 10  5  9  4  9  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 27557.  -3124.  54674.  66459. -13756. -35591.  57622. -65786.], 
        // Q{mac}=[26  0 53 64  0  0 56  0]

        sign=8'b01001111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001001, 8'b00001000, 8'b00001010, 8'b00000101, 8'b00001001, 8'b00000100, 8'b00001001, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001100;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 344: 
        // x=-121, 
        // s=[-1.  1. -1. -1.  1. -1.  1.  1.],
        // w=[ 6  2  3  3 14  3  4  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 28283.  -3366.  55037.  66822. -15450. -35228.  57138. -66391.], 
        // Q{mac}=[27  0 53 65  0  0 55  0]

        sign=8'b01001011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000110, 8'b00000010, 8'b00000011, 8'b00000011, 8'b00001110, 8'b00000011, 8'b00000100, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000111;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 345: 
        // x=-119, 
        // s=[-1.  1.  1. -1.  1. -1.  1.  1.],
        // w=[ 6  3  2 11 10  6  2  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 28997.  -3723.  54799.  68131. -16640. -34514.  56900. -66986.], 
        // Q{mac}=[28  0 53 66  0  0 55  0]

        sign=8'b01101011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000110, 8'b00000011, 8'b00000010, 8'b00001011, 8'b00001010, 8'b00000110, 8'b00000010, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 346: 
        // x=-119, 
        // s=[-1. -1. -1.  1.  1.  1.  1.  1.],
        // w=[4 1 1 3 3 8 5 8],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 29473.  -3604.  54918.  67774. -16997. -35466.  56305. -67938.], 
        // Q{mac}=[28  0 53 66  0  0 54  0]

        sign=8'b00011111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000100, 8'b00000001, 8'b00000001, 8'b00000011, 8'b00000011, 8'b00001000, 8'b00000101, 8'b00001000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 347: 
        // x=-121, 
        // s=[-1. -1.  1.  1.  1.  1. -1.  1.],
        // w=[13 13 13  7 14  3  7 10],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 31046.  -2031.  53345.  66927. -18691. -35829.  57152. -69148.], 
        // Q{mac}=[30  0 52 65  0  0 55  0]

        sign=8'b00111101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001101, 8'b00001101, 8'b00001101, 8'b00000111, 8'b00001110, 8'b00000011, 8'b00000111, 8'b00001010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000111;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 348: 
        // x=-122, 
        // s=[-1. -1. -1.  1.  1.  1.  1. -1.],
        // w=[ 1  6  8  2 10  0  3  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 31168.  -1299.  54321.  66683. -19911. -35829.  56786. -68538.], 
        // Q{mac}=[30  0 53 65  0  0 55  0]

        sign=8'b00011110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00000110, 8'b00001000, 8'b00000010, 8'b00001010, 8'b00000000, 8'b00000011, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 349: 
        // x=-115, 
        // s=[-1. -1. -1. -1.  1.  1.  1.  1.],
        // w=[ 2  5  2  1  5 12  4  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 31398.   -724.  54551.  66798. -20486. -37209.  56326. -68768.], 
        // Q{mac}=[30  0 53 65  0  0 55  0]

        sign=8'b00001111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00000101, 8'b00000010, 8'b00000001, 8'b00000101, 8'b00001100, 8'b00000100, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 350: 
        // x=-121, 
        // s=[-1. -1.  1.  1.  1. -1.  1.  1.],
        // w=[13  8  2  0  8  3  8  7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 32971.    244.  54309.  66798. -21454. -36846.  55358. -69615.], 
        // Q{mac}=[32  0 53 65  0  0 54  0]

        sign=8'b00111011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001101, 8'b00001000, 8'b00000010, 8'b00000000, 8'b00001000, 8'b00000011, 8'b00001000, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000111;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 351: 
        // x=-121, 
        // s=[-1. -1. -1. -1.  1. -1.  1. -1.],
        // w=[ 7  4  7  3 11  9  3  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 33818.    728.  55156.  67161. -22785. -35757.  54995. -69373.], 
        // Q{mac}=[33  0 53 65  0  0 53  0]

        sign=8'b00001010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00000100, 8'b00000111, 8'b00000011, 8'b00001011, 8'b00001001, 8'b00000011, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000111;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 352: 
        // x=-122, 
        // s=[ 1.  1.  1. -1.  1. -1.  1.  1.],
        // w=[0 2 1 4 9 4 5 0],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 33818.    484.  55034.  67649. -23883. -35269.  54385. -69373.], 
        // Q{mac}=[33  0 53 66  0  0 53  0]

        sign=8'b11101011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000000, 8'b00000010, 8'b00000001, 8'b00000100, 8'b00001001, 8'b00000100, 8'b00000101, 8'b00000000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 353: 
        // x=-123, 
        // s=[-1. -1.  1. -1.  1. -1.  1.  1.],
        // w=[ 2  4  0  4 12 13  3  8],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 34064.    976.  55034.  68141. -25359. -33670.  54016. -70357.], 
        // Q{mac}=[33  0 53 66  0  0 52  0]

        sign=8'b00101011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00000100, 8'b00000000, 8'b00000100, 8'b00001100, 8'b00001101, 8'b00000011, 8'b00001000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 354: 
        // x=-123, 
        // s=[ 1. -1.  1. -1. -1. -1. -1.  1.],
        // w=[ 0  5  4  2  1 13  1  4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 34064.   1591.  54542.  68387. -25236. -32071.  54139. -70849.], 
        // Q{mac}=[33  1 53 66  0  0 52  0]

        sign=8'b10100001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000000, 8'b00000101, 8'b00000100, 8'b00000010, 8'b00000001, 8'b00001101, 8'b00000001, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 355: 
        // x=-121, 
        // s=[-1. -1. -1.  1. -1.  1.  1. -1.],
        // w=[3 7 2 3 2 1 3 4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 34427.   2438.  54784.  68024. -24994. -32192.  53776. -70365.], 
        // Q{mac}=[33  2 53 66  0  0 52  0]

        sign=8'b00010110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00000111, 8'b00000010, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000011, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000111;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 356: 
        // x=-127, 
        // s=[ 1. -1.  1. -1.  1.  1. -1. -1.],
        // w=[ 0  3  4  9  0 10  2  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 34427.   2819.  54276.  69167. -24994. -33462.  54030. -69984.], 
        // Q{mac}=[33  2 53 67  0  0 52  0]

        sign=8'b10101100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000000, 8'b00000011, 8'b00000100, 8'b00001001, 8'b00000000, 8'b00001010, 8'b00000010, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 357: 
        // x=-126, 
        // s=[ 1. -1. -1. -1. -1.  1. -1.  1.],
        // w=[0 7 8 1 5 3 1 3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 34427.   3701.  55284.  69293. -24364. -33840.  54156. -70362.], 
        // Q{mac}=[33  3 53 67  0  0 52  0]

        sign=8'b10000101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000000, 8'b00000111, 8'b00001000, 8'b00000001, 8'b00000101, 8'b00000011, 8'b00000001, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 358: 
        // x=-116, 
        // s=[-1.  1. -1. -1.  1.  1.  1.  1.],
        // w=[ 6  5  7  4 15  4  9  0],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 35123.   3121.  56096.  69757. -26104. -34304.  53112. -70362.], 
        // Q{mac}=[34  3 54 68  0  0 51  0]

        sign=8'b01001111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000110, 8'b00000101, 8'b00000111, 8'b00000100, 8'b00001111, 8'b00000100, 8'b00001001, 8'b00000000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001100;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 359: 
        // x=-128, 
        // s=[-1. -1.  1. -1.  1.  1.  1.  1.],
        // w=[1 6 2 1 6 1 6 9],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 35251.   3889.  55840.  69885. -26872. -34432.  52344. -71514.], 
        // Q{mac}=[34  3 54 68  0  0 51  0]

        sign=8'b00101111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00000110, 8'b00000010, 8'b00000001, 8'b00000110, 8'b00000001, 8'b00000110, 8'b00001001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 360: 
        // x=-128, 
        // s=[ 1. -1. -1.  1. -1. -1.  1.  1.],
        // w=[ 3  1  1  5  3 10  1  7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 34867.   4017.  55968.  69245. -26488. -33152.  52216. -72410.], 
        // Q{mac}=[34  3 54 67  0  0 50  0]

        sign=8'b10010011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00000001, 8'b00000001, 8'b00000101, 8'b00000011, 8'b00001010, 8'b00000001, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 361: 
        // x=-128, 
        // s=[ 1.  1. -1. -1.  1.  1. -1.  1.],
        // w=[ 0  1  7  4  3  1 10  1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 34867.   3889.  56864.  69757. -26872. -33280.  53496. -72538.], 
        // Q{mac}=[34  3 55 68  0  0 52  0]

        sign=8'b11001101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000000, 8'b00000001, 8'b00000111, 8'b00000100, 8'b00000011, 8'b00000001, 8'b00001010, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 362: 
        // x=-114, 
        // s=[-1.  1.  1. -1.  1.  1.  1. -1.],
        // w=[ 7  3  0 14  1  5 12  4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 35665.   3547.  56864.  71353. -26986. -33850.  52128. -72082.], 
        // Q{mac}=[34  3 55 69  0  0 50  0]

        sign=8'b01101110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00000011, 8'b00000000, 8'b00001110, 8'b00000001, 8'b00000101, 8'b00001100, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 363: 
        // x=-120, 
        // s=[-1.  1. -1. -1.  1.  1. -1.  1.],
        // w=[12  0  5  1 14  0  2  7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 37105.   3547.  57464.  71473. -28666. -33850.  52368. -72922.], 
        // Q{mac}=[36  3 56 69  0  0 51  0]

        sign=8'b01001101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001100, 8'b00000000, 8'b00000101, 8'b00000001, 8'b00001110, 8'b00000000, 8'b00000010, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 364: 
        // x=-123, 
        // s=[-1.  1. -1.  1.  1. -1.  1.  1.],
        // w=[ 2  0  9  1 14 15  5  9],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 37351.   3547.  58571.  71350. -30388. -32005.  51753. -74029.], 
        // Q{mac}=[36  3 57 69  0  0 50  0]

        sign=8'b01011011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00000000, 8'b00001001, 8'b00000001, 8'b00001110, 8'b00001111, 8'b00000101, 8'b00001001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 365: 
        // x=-61, 
        // s=[-1.  1. -1. -1.  1.  1.  1.  1.],
        // w=[17  6  3 17 11  8 14  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 38388.   3181.  58754.  72387. -31059. -32493.  50899. -74212.], 
        // Q{mac}=[37  3 57 70  0  0 49  0]

        sign=8'b01001111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00010001, 8'b00000110, 8'b00000011, 8'b00010001, 8'b00001011, 8'b00001000, 8'b00001110, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11000011;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 366: 
        // x=-87, 
        // s=[-1.  1.  1. -1.  1.  1.  1. -1.],
        // w=[19  4  7  9 16  6 12  1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 40041.   2833.  58145.  73170. -32451. -33015.  49855. -74125.], 
        // Q{mac}=[39  2 56 71  0  0 48  0]

        sign=8'b01101110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00010011, 8'b00000100, 8'b00000111, 8'b00001001, 8'b00010000, 8'b00000110, 8'b00001100, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10101001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 367: 
        // x=-77, 
        // s=[-1.  1. -1. -1.  1. -1.  1. -1.],
        // w=[ 4  2  4  3 36  2  7  8],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 40349.   2679.  58453.  73401. -35223. -32861.  49316. -73509.], 
        // Q{mac}=[39  2 57 71  0  0 48  0]

        sign=8'b01001010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000100, 8'b00000010, 8'b00000100, 8'b00000011, 8'b00100100, 8'b00000010, 8'b00000111, 8'b00001000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10110011;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 368: 
        // x=-67, 
        // s=[-1. -1.  1.  1.  1. -1. -1.  1.],
        // w=[28 25 17 18  1 18  2  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 42225.   4354.  57314.  72195. -35290. -31655.  49450. -73710.], 
        // Q{mac}=[41  4 55 70  0  0 48  0]

        sign=8'b00111001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00011100, 8'b00011001, 8'b00010001, 8'b00010010, 8'b00000001, 8'b00010010, 8'b00000010, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10111101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 369: 
        // x=9, 
        // s=[-1. -1. -1. -1. -1. -1.  1. -1.],
        // w=[ 6  4 13  2  7  6  3  1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 42171.   4318.  57197.  72177. -35353. -31709.  49477. -73719.], 
        // Q{mac}=[41  4 55 70  0  0 48  0]

        sign=8'b00000010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000110, 8'b00000100, 8'b00001101, 8'b00000010, 8'b00000111, 8'b00000110, 8'b00000011, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00001001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 370: 
        // x=40, 
        // s=[-1. -1. -1.  1.  1. -1.  1. -1.],
        // w=[26  8  2  4 11 22  9  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 41131.   3998.  57117.  72337. -34913. -32589.  49837. -73799.], 
        // Q{mac}=[40  3 55 70  0  0 48  0]

        sign=8'b00011010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00011010, 8'b00001000, 8'b00000010, 8'b00000100, 8'b00001011, 8'b00010110, 8'b00001001, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00101000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 371: 
        // x=57, 
        // s=[ 1. -1. -1.  1. -1. -1.  1. -1.],
        // w=[ 3 16  2 16 22  1 24  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 41302.   3086.  57003.  73249. -36167. -32646.  51205. -73970.], 
        // Q{mac}=[40  3 55 71  0  0 50  0]

        sign=8'b10010010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00010000, 8'b00000010, 8'b00010000, 8'b00010110, 8'b00000001, 8'b00011000, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00111001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 372: 
        // x=16, 
        // s=[-1. -1. -1.  1. -1. -1.  1. -1.],
        // w=[ 2 22  9  3  8  6 17  9],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 41270.   2734.  56859.  73297. -36295. -32742.  51477. -74114.], 
        // Q{mac}=[40  2 55 71  0  0 50  0]

        sign=8'b00010010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00010110, 8'b00001001, 8'b00000011, 8'b00001000, 8'b00000110, 8'b00010001, 8'b00001001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00010000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 373: 
        // x=-24, 
        // s=[-1. -1. -1.  1.  1. -1.  1.  1.],
        // w=[11 13 15  8 19 32 12  4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 41534.   3046.  57219.  73105. -36751. -31974.  51189. -74210.], 
        // Q{mac}=[40  2 55 71  0  0 49  0]

        sign=8'b00011011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001011, 8'b00001101, 8'b00001111, 8'b00001000, 8'b00010011, 8'b00100000, 8'b00001100, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11101000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 374: 
        // x=-75, 
        // s=[ 1.  1.  1. -1.  1. -1. -1. -1.],
        // w=[ 6  4  9  3 22  1 13  4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 41084.   2746.  56544.  73330. -38401. -31899.  52164. -73910.], 
        // Q{mac}=[40  2 55 71  0  0 50  0]

        sign=8'b11101000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000110, 8'b00000100, 8'b00001001, 8'b00000011, 8'b00010110, 8'b00000001, 8'b00001101, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10110101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 375: 
        // x=-117, 
        // s=[ 1.  1. -1. -1.  1. -1. -1.  1.],
        // w=[ 8  3 14 12  3  2  8  1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 40148.   2395.  58182.  74734. -38752. -31665.  53100. -74027.], 
        // Q{mac}=[39  2 56 72  0  0 51  0]

        sign=8'b11001001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001000, 8'b00000011, 8'b00001110, 8'b00001100, 8'b00000011, 8'b00000010, 8'b00001000, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001011;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 376: 
        // x=-81, 
        // s=[ 1. -1.  1. -1.  1. -1. -1.  1.],
        // w=[ 1  2 23  2  9  5 10  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 40067.   2557.  56319.  74896. -39481. -31260.  53910. -74432.], 
        // Q{mac}=[39  2 54 73  0  0 52  0]

        sign=8'b10101001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00000010, 8'b00010111, 8'b00000010, 8'b00001001, 8'b00000101, 8'b00001010, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10101111;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 377: 
        // x=-121, 
        // s=[-1. -1.  1.  1. -1. -1. -1.  1.],
        // w=[2 8 6 7 3 5 5 5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 40309.   3525.  55593.  74049. -39118. -30655.  54515. -75037.], 
        // Q{mac}=[39  3 54 72  0  0 53  0]

        sign=8'b00110001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00001000, 8'b00000110, 8'b00000111, 8'b00000011, 8'b00000101, 8'b00000101, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000111;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 378: 
        // x=-85, 
        // s=[-1. -1.  1.  1.  1.  1. -1. -1.],
        // w=[ 2  2 11  6  4  5 10  1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 40479.   3695.  54658.  73539. -39458. -31080.  55365. -74952.], 
        // Q{mac}=[39  3 53 71  0  0 54  0]

        sign=8'b00111100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00000010, 8'b00001011, 8'b00000110, 8'b00000100, 8'b00000101, 8'b00001010, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10101011;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 379: 
        // x=-117, 
        // s=[ 1. -1.  1. -1. -1. -1. -1.  1.],
        // w=[ 0  1  3  3 12  3  2  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 40479.   3812.  54307.  73890. -38054. -30729.  55599. -75186.], 
        // Q{mac}=[39  3 53 72  0  0 54  0]

        sign=8'b10100001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000000, 8'b00000001, 8'b00000011, 8'b00000011, 8'b00001100, 8'b00000011, 8'b00000010, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001011;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 380: 
        // x=-128, 
        // s=[ 1. -1. -1.  1.  1. -1. -1. -1.],
        // w=[ 3  1 13  1  5  9  4  1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 40095.   3940.  55971.  73762. -38694. -29577.  56111. -75058.], 
        // Q{mac}=[39  3 54 72  0  0 54  0]

        sign=8'b10011000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00000001, 8'b00001101, 8'b00000001, 8'b00000101, 8'b00001001, 8'b00000100, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 381: 
        // x=-128, 
        // s=[-1. -1.  1.  1. -1. -1. -1. -1.],
        // w=[9 8 6 1 1 6 9 5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 41247.   4964.  55203.  73634. -38566. -28809.  57263. -74418.], 
        // Q{mac}=[40  4 53 71  0  0 55  0]

        sign=8'b00110000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001001, 8'b00001000, 8'b00000110, 8'b00000001, 8'b00000001, 8'b00000110, 8'b00001001, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 382: 
        // x=-128, 
        // s=[-1. -1. -1. -1.  1. -1.  1.  1.],
        // w=[3 5 8 2 0 7 7 6],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 41631.   5604.  56227.  73890. -38566. -27913.  56367. -75186.], 
        // Q{mac}=[40  5 54 72  0  0 55  0]

        sign=8'b00001011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00000101, 8'b00001000, 8'b00000010, 8'b00000000, 8'b00000111, 8'b00000111, 8'b00000110};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 383: 
        // x=-128, 
        // s=[ 1.  1.  1. -1. -1. -1. -1. -1.],
        // w=[ 3  2  4  1 10  6  7  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 41247.   5348.  55715.  74018. -37286. -27145.  57263. -74546.], 
        // Q{mac}=[40  5 54 72  0  0 55  0]

        sign=8'b11100000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00000010, 8'b00000100, 8'b00000001, 8'b00001010, 8'b00000110, 8'b00000111, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 384: 
        // x=-128, 
        // s=[-1.  1.  1. -1. -1.  1.  1.  1.],
        // w=[2 7 3 1 6 3 2 1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 41503.   4452.  55331.  74146. -36518. -27529.  57007. -74674.], 
        // Q{mac}=[40  4 54 72  0  0 55  0]

        sign=8'b01100111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00000111, 8'b00000011, 8'b00000001, 8'b00000110, 8'b00000011, 8'b00000010, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 385: 
        // x=-127, 
        // s=[-1. -1. -1. -1. -1. -1.  1.  1.],
        // w=[ 6  1  3 12 11  1  0  7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 42265.   4579.  55712.  75670. -35121. -27402.  57007. -75563.], 
        // Q{mac}=[41  4 54 73  0  0 55  0]

        sign=8'b00000011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000110, 8'b00000001, 8'b00000011, 8'b00001100, 8'b00001011, 8'b00000001, 8'b00000000, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 386: 
        // x=-127, 
        // s=[-1.  1. -1. -1.  1. -1.  1.  1.],
        // w=[ 1  2  9 10  4  1  6  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 42392.   4325.  56855.  76940. -35629. -27275.  56245. -75817.], 
        // Q{mac}=[41  4 55 75  0  0 54  0]

        sign=8'b01001011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00000010, 8'b00001001, 8'b00001010, 8'b00000100, 8'b00000001, 8'b00000110, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 387: 
        // x=-128, 
        // s=[ 1. -1. -1.  1. -1. -1. -1.  1.],
        // w=[1 1 1 0 6 3 8 9],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 42264.   4453.  56983.  76940. -34861. -26891.  57269. -76969.], 
        // Q{mac}=[41  4 55 75  0  0 55  0]

        sign=8'b10010001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00000001, 8'b00000001, 8'b00000000, 8'b00000110, 8'b00000011, 8'b00001000, 8'b00001001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 388: 
        // x=-128, 
        // s=[ 1.  1.  1. -1. -1. -1.  1.  1.],
        // w=[2 3 7 6 2 8 7 7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 42008.   4069.  56087.  77708. -34605. -25867.  56373. -77865.], 
        // Q{mac}=[41  3 54 75  0  0 55  0]

        sign=8'b11100011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00000011, 8'b00000111, 8'b00000110, 8'b00000010, 8'b00001000, 8'b00000111, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 389: 
        // x=-128, 
        // s=[ 1. -1.  1. -1. -1. -1. -1.  1.],
        // w=[0 2 5 8 2 3 3 0],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 42008.   4325.  55447.  78732. -34349. -25483.  56757. -77865.], 
        // Q{mac}=[41  4 54 76  0  0 55  0]

        sign=8'b10100001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000000, 8'b00000010, 8'b00000101, 8'b00001000, 8'b00000010, 8'b00000011, 8'b00000011, 8'b00000000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 390: 
        // x=-127, 
        // s=[ 1.  1. -1. -1.  1. -1. -1.  1.],
        // w=[4 4 9 3 0 1 1 4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 41500.   3817.  56590.  79113. -34349. -25356.  56884. -78373.], 
        // Q{mac}=[40  3 55 77  0  0 55  0]

        sign=8'b11001001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000100, 8'b00000100, 8'b00001001, 8'b00000011, 8'b00000000, 8'b00000001, 8'b00000001, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 391: 
        // x=-127, 
        // s=[-1. -1.  1.  1. -1.  1. -1.  1.],
        // w=[2 4 1 4 8 4 8 9],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 41754.   4325.  56463.  78605. -33333. -25864.  57900. -79516.], 
        // Q{mac}=[40  4 55 76  0  0 56  0]

        sign=8'b00110101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00000100, 8'b00000001, 8'b00000100, 8'b00001000, 8'b00000100, 8'b00001000, 8'b00001001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 392: 
        // x=-128, 
        // s=[ 1.  1. -1.  1.  1. -1.  1. -1.],
        // w=[1 6 5 0 5 9 1 1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 41626.   3557.  57103.  78605. -33973. -24712.  57772. -79388.], 
        // Q{mac}=[40  3 55 76  0  0 56  0]

        sign=8'b11011010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00000110, 8'b00000101, 8'b00000000, 8'b00000101, 8'b00001001, 8'b00000001, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 393: 
        // x=-127, 
        // s=[-1.  1. -1. -1. -1. -1.  1. -1.],
        // w=[ 7  3 11 11  9  1  7  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 42515.   3176.  58500.  80002. -32830. -24585.  56883. -78753.], 
        // Q{mac}=[41  3 57 78  0  0 55  0]

        sign=8'b01000010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00000011, 8'b00001011, 8'b00001011, 8'b00001001, 8'b00000001, 8'b00000111, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 394: 
        // x=-128, 
        // s=[-1.  1. -1. -1. -1.  1. -1.  1.],
        // w=[ 8  2  7  6  9 11  2  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 43539.   2920.  59396.  80770. -31678. -25993.  57139. -79393.], 
        // Q{mac}=[42  2 58 78  0  0 55  0]

        sign=8'b01000101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001000, 8'b00000010, 8'b00000111, 8'b00000110, 8'b00001001, 8'b00001011, 8'b00000010, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 395: 
        // x=-128, 
        // s=[-1. -1.  1.  1. -1.  1. -1.  1.],
        // w=[2 4 0 0 1 1 8 9],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 43795.   3432.  59396.  80770. -31550. -26121.  58163. -80545.], 
        // Q{mac}=[42  3 58 78  0  0 56  0]

        sign=8'b00110101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000001, 8'b00001000, 8'b00001001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 396: 
        // x=-128, 
        // s=[-1. -1.  1.  1. -1. -1. -1.  1.],
        // w=[2 4 4 0 2 4 8 0],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 44051.   3944.  58884.  80770. -31294. -25609.  59187. -80545.], 
        // Q{mac}=[43  3 57 78  0  0 57  0]

        sign=8'b00110001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00000100, 8'b00000100, 8'b00000000, 8'b00000010, 8'b00000100, 8'b00001000, 8'b00000000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 397: 
        // x=-128, 
        // s=[-1.  1. -1.  1. -1. -1. -1.  1.],
        // w=[9 1 2 0 5 9 3 5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 45203.   3816.  59140.  80770. -30654. -24457.  59571. -81185.], 
        // Q{mac}=[44  3 57 78  0  0 58  0]

        sign=8'b01010001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001001, 8'b00000001, 8'b00000010, 8'b00000000, 8'b00000101, 8'b00001001, 8'b00000011, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 398: 
        // x=-128, 
        // s=[-1.  1.  1.  1.  1. -1. -1. -1.],
        // w=[2 4 7 0 0 5 8 5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 45459.   3304.  58244.  80770. -30654. -23817.  60595. -80545.], 
        // Q{mac}=[44  3 56 78  0  0 59  0]

        sign=8'b01111000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00000100, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000101, 8'b00001000, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 399: 
        // x=-128, 
        // s=[ 1.  1.  1.  1.  1.  1. -1.  1.],
        // w=[3 0 3 0 1 3 4 6],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 45075.   3304.  57860.  80770. -30782. -24201.  61107. -81313.], 
        // Q{mac}=[44  3 56 78  0  0 59  0]

        sign=8'b11111101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00000000, 8'b00000011, 8'b00000000, 8'b00000001, 8'b00000011, 8'b00000100, 8'b00000110};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 400: 
        // x=-128, 
        // s=[-1.  1.  1.  1.  1. -1. -1. -1.],
        // w=[9 5 5 7 6 2 3 2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 46227.   2664.  57220.  79874. -31550. -23945.  61491. -81057.], 
        // Q{mac}=[45  2 55 78  0  0 60  0]

        sign=8'b01111000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001001, 8'b00000101, 8'b00000101, 8'b00000111, 8'b00000110, 8'b00000010, 8'b00000011, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 401: 
        // x=-128, 
        // s=[-1. -1. -1.  1. -1. -1. -1.  1.],
        // w=[ 7  4  1  2 12  8  3  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 47123.   3176.  57348.  79618. -30014. -22921.  61875. -81697.], 
        // Q{mac}=[46  3 56 77  0  0 60  0]

        sign=8'b00010001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00000100, 8'b00000001, 8'b00000010, 8'b00001100, 8'b00001000, 8'b00000011, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 402: 
        // x=-128, 
        // s=[-1.  1.  1. -1. -1. -1. -1. -1.],
        // w=[ 8  3 10  3  1 11  2  4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 48147.   2792.  56068.  80002. -29886. -21513.  62131. -81185.], 
        // Q{mac}=[47  2 54 78  0  0 60  0]

        sign=8'b01100000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001000, 8'b00000011, 8'b00001010, 8'b00000011, 8'b00000001, 8'b00001011, 8'b00000010, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 403: 
        // x=-128, 
        // s=[-1.  1. -1. -1. -1.  1. -1.  1.],
        // w=[6 2 2 4 3 1 8 3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 48915.   2536.  56324.  80514. -29502. -21641.  63155. -81569.], 
        // Q{mac}=[47  2 55 78  0  0 61  0]

        sign=8'b01000101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000110, 8'b00000010, 8'b00000010, 8'b00000100, 8'b00000011, 8'b00000001, 8'b00001000, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 404: 
        // x=-128, 
        // s=[ 1. -1. -1.  1. -1. -1. -1.  1.],
        // w=[3 6 8 6 6 8 5 4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 48531.   3304.  57348.  79746. -28734. -20617.  63795. -82081.], 
        // Q{mac}=[47  3 56 77  0  0 62  0]

        sign=8'b10010001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00000110, 8'b00001000, 8'b00000110, 8'b00000110, 8'b00001000, 8'b00000101, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 405: 
        // x=-128, 
        // s=[ 1. -1.  1.  1.  1. -1. -1. -1.],
        // w=[5 8 2 2 5 5 6 2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 47891.   4328.  57092.  79490. -29374. -19977.  64563. -81825.], 
        // Q{mac}=[46  4 55 77  0  0 63  0]

        sign=8'b10111000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000101, 8'b00001000, 8'b00000010, 8'b00000010, 8'b00000101, 8'b00000101, 8'b00000110, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 406: 
        // x=-128, 
        // s=[-1. -1.  1. -1.  1. -1. -1. -1.],
        // w=[9 5 3 2 8 6 2 2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 49043.   4968.  56708.  79746. -30398. -19209.  64819. -81569.], 
        // Q{mac}=[47  4 55 77  0  0 63  0]

        sign=8'b00101000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001001, 8'b00000101, 8'b00000011, 8'b00000010, 8'b00001000, 8'b00000110, 8'b00000010, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 407: 
        // x=-128, 
        // s=[-1.  1. -1.  1. -1. -1. -1.  1.],
        // w=[6 4 3 5 5 9 3 0],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 49811.   4456.  57092.  79106. -29758. -18057.  65203. -81569.], 
        // Q{mac}=[48  4 55 77  0  0 63  0]

        sign=8'b01010001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000110, 8'b00000100, 8'b00000011, 8'b00000101, 8'b00000101, 8'b00001001, 8'b00000011, 8'b00000000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 408: 
        // x=-128, 
        // s=[-1.  1. -1. -1.  1. -1. -1.  1.],
        // w=[4 3 6 7 0 5 5 0],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 50323.   4072.  57860.  80002. -29758. -17417.  65843. -81569.], 
        // Q{mac}=[49  3 56 78  0  0 64  0]

        sign=8'b01001001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000100, 8'b00000011, 8'b00000110, 8'b00000111, 8'b00000000, 8'b00000101, 8'b00000101, 8'b00000000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 409: 
        // x=-128, 
        // s=[-1.  1. -1. -1. -1. -1. -1.  1.],
        // w=[12  5  8  8  9  1  5  9],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 51859.   3432.  58884.  81026. -28606. -17289.  66483. -82721.], 
        // Q{mac}=[50  3 57 79  0  0 64  0]

        sign=8'b01000001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001100, 8'b00000101, 8'b00001000, 8'b00001000, 8'b00001001, 8'b00000001, 8'b00000101, 8'b00001001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 410: 
        // x=-128, 
        // s=[-1. -1. -1.  1.  1. -1.  1.  1.],
        // w=[9 6 7 6 0 7 3 7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 53011.   4200.  59780.  80258. -28606. -16393.  66099. -83617.], 
        // Q{mac}=[51  4 58 78  0  0 64  0]

        sign=8'b00011011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001001, 8'b00000110, 8'b00000111, 8'b00000110, 8'b00000000, 8'b00000111, 8'b00000011, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 411: 
        // x=-128, 
        // s=[ 1.  1. -1. -1.  1. -1. -1. -1.],
        // w=[7 1 1 3 1 4 2 2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 52115.   4072.  59908.  80642. -28734. -15881.  66355. -83361.], 
        // Q{mac}=[50  3 58 78  0  0 64  0]

        sign=8'b11001000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00000001, 8'b00000001, 8'b00000011, 8'b00000001, 8'b00000100, 8'b00000010, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 412: 
        // x=-128, 
        // s=[-1.  1.  1.  1. -1. -1. -1. -1.],
        // w=[4 2 0 3 2 1 6 1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 52627.   3816.  59908.  80258. -28478. -15753.  67123. -83233.], 
        // Q{mac}=[51  3 58 78  0  0 65  0]

        sign=8'b01110000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000100, 8'b00000010, 8'b00000000, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00000110, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 413: 
        // x=-128, 
        // s=[-1.  1.  1.  1. -1.  1.  1. -1.],
        // w=[4 3 1 1 6 0 0 4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 53139.   3432.  59780.  80130. -27710. -15753.  67123. -82721.], 
        // Q{mac}=[51  3 58 78  0  0 65  0]

        sign=8'b01110110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000100, 8'b00000011, 8'b00000001, 8'b00000001, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 414: 
        // x=-128, 
        // s=[-1.  1. -1. -1. -1. -1. -1.  1.],
        // w=[ 1  6  2  2  5 10  6  4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 53267.   2664.  60036.  80386. -27070. -14473.  67891. -83233.], 
        // Q{mac}=[52  2 58 78  0  0 66  0]

        sign=8'b01000001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00000110, 8'b00000010, 8'b00000010, 8'b00000101, 8'b00001010, 8'b00000110, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 415: 
        // x=-128, 
        // s=[-1. -1. -1. -1.  1. -1.  1. -1.],
        // w=[ 6  3  5 11  3  5  5  6],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 54035.   3048.  60676.  81794. -27454. -13833.  67251. -82465.], 
        // Q{mac}=[52  2 59 79  0  0 65  0]

        sign=8'b00001010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000110, 8'b00000011, 8'b00000101, 8'b00001011, 8'b00000011, 8'b00000101, 8'b00000101, 8'b00000110};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 416: 
        // x=-128, 
        // s=[-1. -1.  1.  1.  1. -1. -1.  1.],
        // w=[10  1  3  0  5  8  7  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 55315.   3176.  60292.  81794. -28094. -12809.  68147. -82849.], 
        // Q{mac}=[54  3 58 79  0  0 66  0]

        sign=8'b00111001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001010, 8'b00000001, 8'b00000011, 8'b00000000, 8'b00000101, 8'b00001000, 8'b00000111, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 417: 
        // x=-128, 
        // s=[-1.  1.  1. -1.  1.  1. -1.  1.],
        // w=[2 1 4 2 1 1 8 8],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 55571.   3048.  59780.  82050. -28222. -12937.  69171. -83873.], 
        // Q{mac}=[54  2 58 80  0  0 67  0]

        sign=8'b01101101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00000001, 8'b00000100, 8'b00000010, 8'b00000001, 8'b00000001, 8'b00001000, 8'b00001000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 418: 
        // x=-128, 
        // s=[ 1. -1. -1. -1.  1. -1. -1.  1.],
        // w=[ 1  7  7  5  1  5 10  1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 55443.   3944.  60676.  82690. -28350. -12297.  70451. -84001.], 
        // Q{mac}=[54  3 59 80  0  0 68  0]

        sign=8'b10001001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00000111, 8'b00000111, 8'b00000101, 8'b00000001, 8'b00000101, 8'b00001010, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 419: 
        // x=-128, 
        // s=[-1.  1. -1. -1. -1.  1.  1.  1.],
        // w=[3 6 9 1 4 2 3 2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 55827.   3176.  61828.  82818. -27838. -12553.  70067. -84257.], 
        // Q{mac}=[54  3 60 80  0  0 68  0]

        sign=8'b01000111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00000110, 8'b00001001, 8'b00000001, 8'b00000100, 8'b00000010, 8'b00000011, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 420: 
        // x=-128, 
        // s=[ 1.  1. -1. -1.  1. -1. -1.  1.],
        // w=[ 1  4  9  6  5 11  7  9],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 55699.   2664.  62980.  83586. -28478. -11145.  70963. -85409.], 
        // Q{mac}=[54  2 61 81  0  0 69  0]

        sign=8'b11001001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00000100, 8'b00001001, 8'b00000110, 8'b00000101, 8'b00001011, 8'b00000111, 8'b00001001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 421: 
        // x=-128, 
        // s=[-1.  1. -1. -1. -1. -1.  1.  1.],
        // w=[3 2 2 5 6 4 0 7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 56083.   2408.  63236.  84226. -27710. -10633.  70963. -86305.], 
        // Q{mac}=[54  2 61 82  0  0 69  0]

        sign=8'b01000011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00000010, 8'b00000010, 8'b00000101, 8'b00000110, 8'b00000100, 8'b00000000, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 422: 
        // x=-106, 
        // s=[-1. -1. -1. -1. -1. -1.  1. -1.],
        // w=[ 1 11  6 14  5  3  6  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 56189.   3574.  63872.  85710. -27180. -10315.  70327. -86093.], 
        // Q{mac}=[54  3 62 83  0  0 68  0]

        sign=8'b00000010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00001011, 8'b00000110, 8'b00001110, 8'b00000101, 8'b00000011, 8'b00000110, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10010110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 423: 
        // x=-104, 
        // s=[-1.  1.  1. -1.  1. -1. -1. -1.],
        // w=[10  3  3  8 10  4  2  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 57229.   3262.  63560.  86542. -28220.  -9899.  70535. -85573.], 
        // Q{mac}=[55  3 62 84  0  0 68  0]

        sign=8'b01101000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001010, 8'b00000011, 8'b00000011, 8'b00001000, 8'b00001010, 8'b00000100, 8'b00000010, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10011000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 424: 
        // x=-118, 
        // s=[-1.  1. -1. -1. -1.  1.  1. -1.],
        // w=[11  8  5  5  3  4  8  4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 58527.   2318.  64150.  87132. -27866. -10371.  69591. -85101.], 
        // Q{mac}=[57  2 62 85  0  0 67  0]

        sign=8'b01000110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001011, 8'b00001000, 8'b00000101, 8'b00000101, 8'b00000011, 8'b00000100, 8'b00001000, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 425: 
        // x=-116, 
        // s=[-1. -1. -1. -1.  1. -1.  1.  1.],
        // w=[ 7  2  5 15 10  9  0  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 59339.   2550.  64730.  88872. -29026.  -9327.  69591. -85681.], 
        // Q{mac}=[57  2 63 86  0  0 67  0]

        sign=8'b00001011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00000010, 8'b00000101, 8'b00001111, 8'b00001010, 8'b00001001, 8'b00000000, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001100;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 426: 
        // x=-106, 
        // s=[-1. -1.  1.  1. -1.  1.  1.  1.],
        // w=[10  5 13  0  1  1  5  6],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 60399.   3080.  63352.  88872. -28920.  -9433.  69061. -86317.], 
        // Q{mac}=[58  3 61 86  0  0 67  0]

        sign=8'b00110111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001010, 8'b00000101, 8'b00001101, 8'b00000000, 8'b00000001, 8'b00000001, 8'b00000101, 8'b00000110};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10010110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 427: 
        // x=-123, 
        // s=[-1. -1.  1.  1. -1.  1.  1.  1.],
        // w=[13  9  3  3  9  9  6  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 61998.   4187.  62983.  88503. -27813. -10540.  68323. -86932.], 
        // Q{mac}=[60  4 61 86  0  0 66  0]

        sign=8'b00110111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001101, 8'b00001001, 8'b00000011, 8'b00000011, 8'b00001001, 8'b00001001, 8'b00000110, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 428: 
        // x=-111, 
        // s=[ 1. -1. -1. -1.  1.  1.  1.  1.],
        // w=[6 9 1 5 7 5 4 5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 61332.   5186.  63094.  89058. -28590. -11095.  67879. -87487.], 
        // Q{mac}=[59  5 61 86  0  0 66  0]

        sign=8'b10001111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000110, 8'b00001001, 8'b00000001, 8'b00000101, 8'b00000111, 8'b00000101, 8'b00000100, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10010001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 429: 
        // x=-107, 
        // s=[-1.  1.  1.  1.  1. -1.  1. -1.],
        // w=[15  0  2  7  1  6  5  6],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 62937.   5186.  62880.  88309. -28697. -10453.  67344. -86845.], 
        // Q{mac}=[61  5 61 86  0  0 65  0]

        sign=8'b01111010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001111, 8'b00000000, 8'b00000010, 8'b00000111, 8'b00000001, 8'b00000110, 8'b00000101, 8'b00000110};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10010101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 430: 
        // x=-121, 
        // s=[-1. -1. -1. -1.  1.  1. -1.  1.],
        // w=[ 1  5  3  6 14  9  5  0],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 63058.   5791.  63243.  89035. -30391. -11542.  67949. -86845.], 
        // Q{mac}=[61  5 61 86  0  0 66  0]

        sign=8'b00001101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00000101, 8'b00000011, 8'b00000110, 8'b00001110, 8'b00001001, 8'b00000101, 8'b00000000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000111;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 431: 
        // x=-116, 
        // s=[-1.  1. -1. -1.  1. -1.  1.  1.],
        // w=[ 7  4  7 10 14 10  7  6],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 63870.   5327.  64055.  90195. -32015. -10382.  67137. -87541.], 
        // Q{mac}=[62  5 62 88  0  0 65  0]

        sign=8'b01001011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00000100, 8'b00000111, 8'b00001010, 8'b00001110, 8'b00001010, 8'b00000111, 8'b00000110};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001100;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 432: 
        // x=-113, 
        // s=[-1. -1.  1.  1. -1.  1. -1. -1.],
        // w=[ 7 11  7 11  8  7  6  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 64661.   6570.  63264.  88952. -31111. -11173.  67815. -86976.], 
        // Q{mac}=[63  6 61 86  0  0 66  0]

        sign=8'b00110100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00001011, 8'b00000111, 8'b00001011, 8'b00001000, 8'b00000111, 8'b00000110, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001111;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 433: 
        // x=-124, 
        // s=[-1.  1.  1. -1. -1.  1. -1.  1.],
        // w=[13  0  9  4 12 14  1  7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 66273.   6570.  62148.  89448. -29623. -12909.  67939. -87844.], 
        // Q{mac}=[64  6 60 87  0  0 66  0]

        sign=8'b01100101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001101, 8'b00000000, 8'b00001001, 8'b00000100, 8'b00001100, 8'b00001110, 8'b00000001, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000100;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 434: 
        // x=-113, 
        // s=[-1. -1.  1. -1.  1.  1.  1.  1.],
        // w=[2 6 6 6 2 2 4 6],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 66499.   7248.  61470.  90126. -29849. -13135.  67487. -88522.], 
        // Q{mac}=[64  7 60 88  0  0 65  0]

        sign=8'b00101111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00000110, 8'b00000110, 8'b00000110, 8'b00000010, 8'b00000010, 8'b00000100, 8'b00000110};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001111;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 435: 
        // x=-122, 
        // s=[-1.  1.  1.  1. -1.  1. -1. -1.],
        // w=[5 3 4 0 1 5 3 3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 67109.   6882.  60982.  90126. -29727. -13745.  67853. -88156.], 
        // Q{mac}=[65  6 59 88  0  0 66  0]

        sign=8'b01110100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000101, 8'b00000011, 8'b00000100, 8'b00000000, 8'b00000001, 8'b00000101, 8'b00000011, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 436: 
        // x=-118, 
        // s=[ 1. -1.  1.  1. -1.  1. -1.  1.],
        // w=[4 3 3 3 6 9 9 4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 66637.   7236.  60628.  89772. -29019. -14807.  68915. -88628.], 
        // Q{mac}=[65  7 59 87  0  0 67  0]

        sign=8'b10110101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000100, 8'b00000011, 8'b00000011, 8'b00000011, 8'b00000110, 8'b00001001, 8'b00001001, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 437: 
        // x=-107, 
        // s=[-1. -1.  1. -1.  1.  1.  1.  1.],
        // w=[7 6 3 8 3 9 1 0],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 67386.   7878.  60307.  90628. -29340. -15770.  68808. -88628.], 
        // Q{mac}=[65  7 58 88  0  0 67  0]

        sign=8'b00101111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00000110, 8'b00000011, 8'b00001000, 8'b00000011, 8'b00001001, 8'b00000001, 8'b00000000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10010101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 438: 
        // x=-128, 
        // s=[-1. -1. -1. -1.  1.  1.  1.  1.],
        // w=[3 4 5 8 0 2 5 2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 67770.   8390.  60947.  91652. -29340. -16026.  68168. -88884.], 
        // Q{mac}=[66  8 59 89  0  0 66  0]

        sign=8'b00001111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00000100, 8'b00000101, 8'b00001000, 8'b00000000, 8'b00000010, 8'b00000101, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 439: 
        // x=-126, 
        // s=[-1.  1.  1.  1. -1. -1. -1.  1.],
        // w=[7 3 2 7 5 3 5 0],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 68652.   8012.  60695.  90770. -28710. -15648.  68798. -88884.], 
        // Q{mac}=[67  7 59 88  0  0 67  0]

        sign=8'b01110001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00000011, 8'b00000010, 8'b00000111, 8'b00000101, 8'b00000011, 8'b00000101, 8'b00000000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 440: 
        // x=-128, 
        // s=[-1.  1.  1. -1. -1.  1.  1.  1.],
        // w=[11  5  8  1  9  2  0  8],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 70060.   7372.  59671.  90898. -27558. -15904.  68798. -89908.], 
        // Q{mac}=[68  7 58 88  0  0 67  0]

        sign=8'b01100111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001011, 8'b00000101, 8'b00001000, 8'b00000001, 8'b00001001, 8'b00000010, 8'b00000000, 8'b00001000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 441: 
        // x=-113, 
        // s=[ 1. -1.  1. -1. -1.  1.  1.  1.],
        // w=[ 0  9  7  7  9 20  6  7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 70060.   8389.  58880.  91689. -26541. -18164.  68120. -90699.], 
        // Q{mac}=[68  8 57 89  0  0 66  0]

        sign=8'b10100111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000000, 8'b00001001, 8'b00000111, 8'b00000111, 8'b00001001, 8'b00010100, 8'b00000110, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001111;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 442: 
        // x=-108, 
        // s=[-1.  1.  1. -1. -1.  1. -1.  1.],
        // w=[9 7 1 3 2 4 5 7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 71032.   7633.  58772.  92013. -26325. -18596.  68660. -91455.], 
        // Q{mac}=[69  7 57 89  0  0 67  0]

        sign=8'b01100101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001001, 8'b00000111, 8'b00000001, 8'b00000011, 8'b00000010, 8'b00000100, 8'b00000101, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10010100;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 443: 
        // x=-119, 
        // s=[ 1.  1. -1. -1. -1.  1.  1.  1.],
        // w=[ 2  8  8 10 13  7  9  0],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 70794.   6681.  59724.  93203. -24778. -19429.  67589. -91455.], 
        // Q{mac}=[69  6 58 91  0  0 66  0]

        sign=8'b11000111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00001000, 8'b00001000, 8'b00001010, 8'b00001101, 8'b00000111, 8'b00001001, 8'b00000000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 444: 
        // x=-1, 
        // s=[-1. -1. -1.  1.  1.  1.  1. -1.],
        // w=[18 33 20 12  3 10 37  1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 70812.   6714.  59744.  93191. -24781. -19439.  67552. -91454.], 
        // Q{mac}=[69  6 58 91  0  0 65  0]

        sign=8'b00011110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00010010, 8'b00100001, 8'b00010100, 8'b00001100, 8'b00000011, 8'b00001010, 8'b00100101, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11111111;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 445: 
        // x=25, 
        // s=[ 1.  1. -1. -1.  1.  1. -1.  1.],
        // w=[ 7 12  2  2 13 10  7  0],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 70987.   7014.  59694.  93141. -24456. -19189.  67377. -91454.], 
        // Q{mac}=[69  6 58 90  0  0 65  0]

        sign=8'b11001101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00001100, 8'b00000010, 8'b00000010, 8'b00001101, 8'b00001010, 8'b00000111, 8'b00000000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00011001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 446: 
        // x=-33, 
        // s=[ 1.  1.  1. -1.  1.  1. -1. -1.],
        // w=[ 0  2  5  5  3 13  2  4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 70987.   6948.  59529.  93306. -24555. -19618.  67443. -91322.], 
        // Q{mac}=[69  6 58 91  0  0 65  0]

        sign=8'b11101100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000000, 8'b00000010, 8'b00000101, 8'b00000101, 8'b00000011, 8'b00001101, 8'b00000010, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11011111;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 447: 
        // x=-128, 
        // s=[ 1. -1.  1.  1. -1. -1. -1. -1.],
        // w=[ 8  8  5  1  4 10  7  1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 69963.   7972.  58889.  93178. -24043. -18338.  68339. -91194.], 
        // Q{mac}=[68  7 57 90  0  0 66  0]

        sign=8'b10110000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001000, 8'b00001000, 8'b00000101, 8'b00000001, 8'b00000100, 8'b00001010, 8'b00000111, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 448: 
        // x=-120, 
        // s=[-1. -1. -1.  1.  1. -1. -1. -1.],
        // w=[12 15  3  5  7 16  2  1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 71403.   9772.  59249.  92578. -24883. -16418.  68579. -91074.], 
        // Q{mac}=[69  9 57 90  0  0 66  0]

        sign=8'b00011000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001100, 8'b00001111, 8'b00000011, 8'b00000101, 8'b00000111, 8'b00010000, 8'b00000010, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 449: 
        // x=-120, 
        // s=[-1. -1.  1.  1.  1. -1. -1. -1.],
        // w=[ 9  4  3 14 17 28  6  1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 72483.  10252.  58889.  90898. -26923. -13058.  69299. -90954.], 
        // Q{mac}=[70 10 57 88  0  0 67  0]

        sign=8'b00111000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001001, 8'b00000100, 8'b00000011, 8'b00001110, 8'b00010001, 8'b00011100, 8'b00000110, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 450: 
        // x=22, 
        // s=[ 1.  1.  1. -1. -1.  1. -1.  1.],
        // w=[ 46  58  43   3  15  17 106   0],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 73495.  11528.  59835.  90832. -27253. -12684.  66967. -90954.], 
        // Q{mac}=[71 11 58 88  0  0 65  0]

        sign=8'b11100101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00101110, 8'b00111010, 8'b00101011, 8'b00000011, 8'b00001111, 8'b00010001, 8'b01101010, 8'b00000000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00010110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 451: 
        // x=-9, 
        // s=[-1. -1. -1.  1. -1.  1.  1.  1.],
        // w=[ 8 19 31 28  9  2 24  7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 73567.  11699.  60114.  90580. -27172. -12702.  66751. -91017.], 
        // Q{mac}=[71 11 58 88  0  0 65  0]

        sign=8'b00010111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001000, 8'b00010011, 8'b00011111, 8'b00011100, 8'b00001001, 8'b00000010, 8'b00011000, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11110111;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 452: 
        // x=55, 
        // s=[ 1.  1. -1.  1.  1. -1. -1. -1.],
        // w=[27 16 19 15 14  4 16  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 75052.  12579.  59069.  91405. -26402. -12922.  65871. -91127.], 
        // Q{mac}=[73 12 57 89  0  0 64  0]

        sign=8'b11011000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00011011, 8'b00010000, 8'b00010011, 8'b00001111, 8'b00001110, 8'b00000100, 8'b00010000, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00110111;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 453: 
        // x=-51, 
        // s=[-1. -1. -1.  1.  1.  1.  1.  1.],
        // w=[ 3  3 27 12  6  0 26  0],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 75205.  12732.  60446.  90793. -26708. -12922.  64545. -91127.], 
        // Q{mac}=[73 12 59 88  0  0 63  0]

        sign=8'b00011111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00000011, 8'b00011011, 8'b00001100, 8'b00000110, 8'b00000000, 8'b00011010, 8'b00000000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11001101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 454: 
        // x=-90, 
        // s=[-1.  1. -1. -1. -1.  1.  1.  1.],
        // w=[ 1  9 16  4  3  7  8  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 75295.  11922.  61886.  91153. -26438. -13552.  63825. -91577.], 
        // Q{mac}=[73 11 60 89  0  0 62  0]

        sign=8'b01000111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00001001, 8'b00010000, 8'b00000100, 8'b00000011, 8'b00000111, 8'b00001000, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10100110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 455: 
        // x=-50, 
        // s=[ 1.  1.  1.  1. -1.  1. -1. -1.],
        // w=[ 6  4 19  7 13 28 24  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 74995.  11722.  60936.  90803. -25788. -14952.  65025. -91327.], 
        // Q{mac}=[73 11 59 88  0  0 63  0]

        sign=8'b11110100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000110, 8'b00000100, 8'b00010011, 8'b00000111, 8'b00001101, 8'b00011100, 8'b00011000, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11001110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 456: 
        // x=-101, 
        // s=[ 1. -1.  1. -1. -1.  1. -1.  1.],
        // w=[ 5  4  4  3 21 21  3  6],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 74490.  12126.  60532.  91106. -23667. -17073.  65328. -91933.], 
        // Q{mac}=[72 11 59 88  0  0 63  0]

        sign=8'b10100101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000101, 8'b00000100, 8'b00000100, 8'b00000011, 8'b00010101, 8'b00010101, 8'b00000011, 8'b00000110};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10011011;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 457: 
        // x=-63, 
        // s=[-1. -1.  1.  1. -1.  1. -1.  1.],
        // w=[ 1 18 37  8 39 46 25  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 74553.  13260.  58201.  90602. -21210. -19971.  66903. -92248.], 
        // Q{mac}=[72 12 56 88  0  0 65  0]

        sign=8'b00110101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00010010, 8'b00100101, 8'b00001000, 8'b00100111, 8'b00101110, 8'b00011001, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11000001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 458: 
        // x=-101, 
        // s=[ 1. -1.  1. -1. -1.  1. -1. -1.],
        // w=[ 3  4 20  4 31 24 18  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 74250.  13664.  56181.  91006. -18079. -22395.  68721. -91945.], 
        // Q{mac}=[72 13 54 88  0  0 67  0]

        sign=8'b10100100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00000100, 8'b00010100, 8'b00000100, 8'b00011111, 8'b00011000, 8'b00010010, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10011011;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 459: 
        // x=-128, 
        // s=[ 1.  1.  1. -1. -1.  1. -1.  1.],
        // w=[9 1 1 5 3 3 4 4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 73098.  13536.  56053.  91646. -17695. -22779.  69233. -92457.], 
        // Q{mac}=[71 13 54 89  0  0 67  0]

        sign=8'b11100101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001001, 8'b00000001, 8'b00000001, 8'b00000101, 8'b00000011, 8'b00000011, 8'b00000100, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 460: 
        // x=-127, 
        // s=[ 1. -1.  1.  1. -1. -1. -1.  1.],
        // w=[ 4 16 12  4  2  4 11  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 72590.  15568.  54529.  91138. -17441. -22271.  70630. -92838.], 
        // Q{mac}=[70 15 53 89  0  0 68  0]

        sign=8'b10110001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000100, 8'b00010000, 8'b00001100, 8'b00000100, 8'b00000010, 8'b00000100, 8'b00001011, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 461: 
        // x=-128, 
        // s=[ 1. -1.  1.  1. -1.  1. -1. -1.],
        // w=[ 5 13  5  4  4  0  8  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 71950.  17232.  53889.  90626. -16929. -22271.  71654. -92582.], 
        // Q{mac}=[70 16 52 88  0  0 69  0]

        sign=8'b10110100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000101, 8'b00001101, 8'b00000101, 8'b00000100, 8'b00000100, 8'b00000000, 8'b00001000, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 462: 
        // x=-128, 
        // s=[-1. -1.  1. -1. -1. -1. -1.  1.],
        // w=[1 2 2 8 2 8 9 6],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 72078.  17488.  53633.  91650. -16673. -21247.  72806. -93350.], 
        // Q{mac}=[70 17 52 89  0  0 71  0]

        sign=8'b00100001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00000010, 8'b00000010, 8'b00001000, 8'b00000010, 8'b00001000, 8'b00001001, 8'b00000110};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 463: 
        // x=-127, 
        // s=[-1.  1.  1. -1. -1. -1. -1.  1.],
        // w=[ 5  1  7  3 11  5  5  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 72713.  17361.  52744.  92031. -15276. -20612.  73441. -93731.], 
        // Q{mac}=[71 16 51 89  0  0 71  0]

        sign=8'b01100001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000101, 8'b00000001, 8'b00000111, 8'b00000011, 8'b00001011, 8'b00000101, 8'b00000101, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 464: 
        // x=-127, 
        // s=[ 1. -1.  1.  1.  1. -1. -1.  1.],
        // w=[ 1  2  2  4  4  1 11  7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 72586.  17615.  52490.  91523. -15784. -20485.  74838. -94620.], 
        // Q{mac}=[70 17 51 89  0  0 73  0]

        sign=8'b10111001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00000010, 8'b00000010, 8'b00000100, 8'b00000100, 8'b00000001, 8'b00001011, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 465: 
        // x=-126, 
        // s=[ 1. -1. -1.  1.  1.  1.  1.  1.],
        // w=[ 1 10  4  5  3  2  1  8],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 72460.  18875.  52994.  90893. -16162. -20737.  74712. -95628.], 
        // Q{mac}=[70 18 51 88  0  0 72  0]

        sign=8'b10011111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00001010, 8'b00000100, 8'b00000101, 8'b00000011, 8'b00000010, 8'b00000001, 8'b00001000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 466: 
        // x=-127, 
        // s=[-1. -1.  1.  1. -1. -1.  1.  1.],
        // w=[3 9 0 1 7 8 3 0],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 72841.  20018.  52994.  90766. -15273. -19721.  74331. -95628.], 
        // Q{mac}=[71 19 51 88  0  0 72  0]

        sign=8'b00110011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00001001, 8'b00000000, 8'b00000001, 8'b00000111, 8'b00001000, 8'b00000011, 8'b00000000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 467: 
        // x=-128, 
        // s=[ 1.  1.  1. -1.  1. -1.  1.  1.],
        // w=[ 8  4  5  6  4 10  4  1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 71817.  19506.  52354.  91534. -15785. -18441.  73819. -95756.], 
        // Q{mac}=[70 19 51 89  0  0 72  0]

        sign=8'b11101011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001000, 8'b00000100, 8'b00000101, 8'b00000110, 8'b00000100, 8'b00001010, 8'b00000100, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 468: 
        // x=-128, 
        // s=[ 1. -1.  1.  1. -1.  1. -1.  1.],
        // w=[ 6  1 11  5 10  6  5  1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 71049.  19634.  50946.  90894. -14505. -19209.  74459. -95884.], 
        // Q{mac}=[69 19 49 88  0  0 72  0]

        sign=8'b10110101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000110, 8'b00000001, 8'b00001011, 8'b00000101, 8'b00001010, 8'b00000110, 8'b00000101, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 469: 
        // x=-127, 
        // s=[ 1. -1.  1.  1.  1. -1.  1. -1.],
        // w=[5 4 1 4 0 4 3 2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 70414.  20142.  50819.  90386. -14505. -18701.  74078. -95630.], 
        // Q{mac}=[68 19 49 88  0  0 72  0]

        sign=8'b10111010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000101, 8'b00000100, 8'b00000001, 8'b00000100, 8'b00000000, 8'b00000100, 8'b00000011, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 470: 
        // x=-127, 
        // s=[ 1. -1.  1.  1. -1. -1.  1.  1.],
        // w=[ 6 10  0  2  8  7  4  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 69652.  21412.  50819.  90132. -13489. -17812.  73570. -96011.], 
        // Q{mac}=[68 20 49 88  0  0 71  0]

        sign=8'b10110011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000110, 8'b00001010, 8'b00000000, 8'b00000010, 8'b00001000, 8'b00000111, 8'b00000100, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 471: 
        // x=-128, 
        // s=[ 1.  1.  1. -1.  1.  1. -1.  1.],
        // w=[ 6  0  2 10  5  4  4  7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 68884.  21412.  50563.  91412. -14129. -18324.  74082. -96907.], 
        // Q{mac}=[67 20 49 89  0  0 72  0]

        sign=8'b11101101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000110, 8'b00000000, 8'b00000010, 8'b00001010, 8'b00000101, 8'b00000100, 8'b00000100, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 472: 
        // x=-128, 
        // s=[ 1. -1.  1. -1. -1.  1.  1. -1.],
        // w=[7 5 5 8 7 3 3 6],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 67988.  22052.  49923.  92436. -13233. -18708.  73698. -96139.], 
        // Q{mac}=[66 21 48 90  0  0 71  0]

        sign=8'b10100110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00000101, 8'b00000101, 8'b00001000, 8'b00000111, 8'b00000011, 8'b00000011, 8'b00000110};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 473: 
        // x=-126, 
        // s=[-1. -1.  1.  1. -1.  1. -1. -1.],
        // w=[12  7 10  3  3  1  4  7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 69500.  22934.  48663.  92058. -12855. -18834.  74202. -95257.], 
        // Q{mac}=[67 22 47 89  0  0 72  0]

        sign=8'b00110100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001100, 8'b00000111, 8'b00001010, 8'b00000011, 8'b00000011, 8'b00000001, 8'b00000100, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 474: 
        // x=-128, 
        // s=[-1.  1.  1.  1.  1.  1. -1.  1.],
        // w=[6 6 6 2 1 3 9 3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 70268.  22166.  47895.  91802. -12983. -19218.  75354. -95641.], 
        // Q{mac}=[68 21 46 89  0  0 73  0]

        sign=8'b01111101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000110, 8'b00000110, 8'b00000110, 8'b00000010, 8'b00000001, 8'b00000011, 8'b00001001, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 475: 
        // x=-128, 
        // s=[-1. -1. -1.  1.  1. -1. -1.  1.],
        // w=[2 1 2 3 4 6 3 8],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 70524.  22294.  48151.  91418. -13495. -18450.  75738. -96665.], 
        // Q{mac}=[68 21 47 89  0  0 73  0]

        sign=8'b00011001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00000001, 8'b00000010, 8'b00000011, 8'b00000100, 8'b00000110, 8'b00000011, 8'b00001000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 476: 
        // x=-128, 
        // s=[ 1.  1. -1. -1. -1.  1. -1.  1.],
        // w=[ 1  7  4 10 10  4  5  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 70396.  21398.  48663.  92698. -12215. -18962.  76378. -97305.], 
        // Q{mac}=[68 20 47 90  0  0 74  0]

        sign=8'b11000101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00000111, 8'b00000100, 8'b00001010, 8'b00001010, 8'b00000100, 8'b00000101, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 477: 
        // x=-128, 
        // s=[-1. -1. -1. -1. -1.  1. -1.  1.],
        // w=[6 4 5 1 5 6 2 4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 71164.  21910.  49303.  92826. -11575. -19730.  76634. -97817.], 
        // Q{mac}=[69 21 48 90  0  0 74  0]

        sign=8'b00000101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000110, 8'b00000100, 8'b00000101, 8'b00000001, 8'b00000101, 8'b00000110, 8'b00000010, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 478: 
        // x=-127, 
        // s=[-1. -1. -1. -1.  1. -1. -1.  1.],
        // w=[ 4  7  1 10  4  9  7  4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 71672.  22799.  49430.  94096. -12083. -18587.  77523. -98325.], 
        // Q{mac}=[69 22 48 91  0  0 75  0]

        sign=8'b00001001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000100, 8'b00000111, 8'b00000001, 8'b00001010, 8'b00000100, 8'b00001001, 8'b00000111, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 479: 
        // x=-127, 
        // s=[-1.  1. -1.  1. -1.  1. -1. -1.],
        // w=[4 1 6 0 8 2 4 3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 72180.  22672.  50192.  94096. -11067. -18841.  78031. -97944.], 
        // Q{mac}=[70 22 49 91  0  0 76  0]

        sign=8'b01010100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000100, 8'b00000001, 8'b00000110, 8'b00000000, 8'b00001000, 8'b00000010, 8'b00000100, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 480: 
        // x=-127, 
        // s=[ 1. -1.  1. -1.  1.  1.  1. -1.],
        // w=[ 0  5  7 10  2  8  6  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 72180.  23307.  49303.  95366. -11321. -19857.  77269. -97563.], 
        // Q{mac}=[70 22 48 93  0  0 75  0]

        sign=8'b10101110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000000, 8'b00000101, 8'b00000111, 8'b00001010, 8'b00000010, 8'b00001000, 8'b00000110, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 481: 
        // x=-126, 
        // s=[-1. -1. -1. -1.  1. -1.  1. -1.],
        // w=[ 4 10  1  5  3  2  3  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 72684.  24567.  49429.  95996. -11699. -19605.  76891. -97185.], 
        // Q{mac}=[70 23 48 93  0  0 75  0]

        sign=8'b00001010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000100, 8'b00001010, 8'b00000001, 8'b00000101, 8'b00000011, 8'b00000010, 8'b00000011, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 482: 
        // x=-128, 
        // s=[-1.  1. -1. -1.  1.  1. -1.  1.],
        // w=[8 3 4 1 3 5 7 8],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 73708.  24183.  49941.  96124. -12083. -20245.  77787. -98209.], 
        // Q{mac}=[71 23 48 93  0  0 75  0]

        sign=8'b01001101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001000, 8'b00000011, 8'b00000100, 8'b00000001, 8'b00000011, 8'b00000101, 8'b00000111, 8'b00001000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 483: 
        // x=-127, 
        // s=[ 1. -1.  1. -1. -1. -1. -1.  1.],
        // w=[5 3 6 1 9 3 1 4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 73073.  24564.  49179.  96251. -10940. -19864.  77914. -98717.], 
        // Q{mac}=[71 23 48 93  0  0 76  0]

        sign=8'b10100001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000101, 8'b00000011, 8'b00000110, 8'b00000001, 8'b00001001, 8'b00000011, 8'b00000001, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 484: 
        // x=-127, 
        // s=[-1. -1. -1. -1. -1. -1. -1.  1.],
        // w=[ 6  1  4  1 11  6  2  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 73835.  24691.  49687.  96378.  -9543. -19102.  78168. -99352.], 
        // Q{mac}=[72 24 48 94  0  0 76  0]

        sign=8'b00000001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000110, 8'b00000001, 8'b00000100, 8'b00000001, 8'b00001011, 8'b00000110, 8'b00000010, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 485: 
        // x=-126, 
        // s=[-1.  1. -1. -1.  1. -1. -1.  1.],
        // w=[13  0  3  6  5 10  7  8],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  75473.   24691.   50065.   97134.  -10173.  -17842.   79050. -100360.], 
        // Q{mac}=[73 24 48 94  0  0 77  0]

        sign=8'b01001001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001101, 8'b00000000, 8'b00000011, 8'b00000110, 8'b00000101, 8'b00001010, 8'b00000111, 8'b00001000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 486: 
        // x=-128, 
        // s=[ 1.  1.  1. -1. -1. -1.  1.  1.],
        // w=[0 7 3 5 6 1 5 1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  75473.   23795.   49681.   97774.   -9405.  -17714.   78410. -100488.], 
        // Q{mac}=[73 23 48 95  0  0 76  0]

        sign=8'b11100011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000000, 8'b00000111, 8'b00000011, 8'b00000101, 8'b00000110, 8'b00000001, 8'b00000101, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 487: 
        // x=-128, 
        // s=[-1. -1.  1.  1. -1.  1.  1. -1.],
        // w=[ 7 12  5  4  9  3  3  7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 76369.  25331.  49041.  97262.  -8253. -18098.  78026. -99592.], 
        // Q{mac}=[74 24 47 94  0  0 76  0]

        sign=8'b00110110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00001100, 8'b00000101, 8'b00000100, 8'b00001001, 8'b00000011, 8'b00000011, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 488: 
        // x=-128, 
        // s=[-1.  1. -1.  1.  1. -1. -1.  1.],
        // w=[2 7 7 1 6 8 1 4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  76625.   24435.   49937.   97134.   -9021.  -17074.   78154. -100104.], 
        // Q{mac}=[74 23 48 94  0  0 76  0]

        sign=8'b01011001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00000111, 8'b00000111, 8'b00000001, 8'b00000110, 8'b00001000, 8'b00000001, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 489: 
        // x=-128, 
        // s=[-1. -1. -1. -1. -1.  1. -1.  1.],
        // w=[ 2  5  7  1 14  4  4  7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  76881.   25075.   50833.   97262.   -7229.  -17586.   78666. -101000.], 
        // Q{mac}=[75 24 49 94  0  0 76  0]

        sign=8'b00000101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00000101, 8'b00000111, 8'b00000001, 8'b00001110, 8'b00000100, 8'b00000100, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 490: 
        // x=-128, 
        // s=[-1. -1. -1. -1. -1. -1. -1. -1.],
        // w=[1 3 5 2 3 9 6 2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  77009.   25459.   51473.   97518.   -6845.  -16434.   79434. -100744.], 
        // Q{mac}=[75 24 50 95  0  0 77  0]

        sign=8'b00000000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000011, 8'b00001001, 8'b00000110, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 491: 
        // x=-128, 
        // s=[-1.  1.  1. -1. -1. -1.  1.  1.],
        // w=[7 6 1 3 8 6 5 9],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  77905.   24691.   51345.   97902.   -5821.  -15666.   78794. -101896.], 
        // Q{mac}=[76 24 50 95  0  0 76  0]

        sign=8'b01100011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00000110, 8'b00000001, 8'b00000011, 8'b00001000, 8'b00000110, 8'b00000101, 8'b00001001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 492: 
        // x=-128, 
        // s=[ 1.  1.  1.  1. -1. -1. -1. -1.],
        // w=[6 4 6 4 5 5 7 2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  77137.   24179.   50577.   97390.   -5181.  -15026.   79690. -101640.], 
        // Q{mac}=[75 23 49 95  0  0 77  0]

        sign=8'b11110000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000110, 8'b00000100, 8'b00000110, 8'b00000100, 8'b00000101, 8'b00000101, 8'b00000111, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 493: 
        // x=-128, 
        // s=[-1. -1.  1.  1. -1. -1. -1. -1.],
        // w=[5 6 4 2 7 2 1 7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  77777.   24947.   50065.   97134.   -4285.  -14770.   79818. -100744.], 
        // Q{mac}=[75 24 48 94  0  0 77  0]

        sign=8'b00110000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000101, 8'b00000110, 8'b00000100, 8'b00000010, 8'b00000111, 8'b00000010, 8'b00000001, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 494: 
        // x=-128, 
        // s=[-1.  1. -1. -1.  1. -1. -1. -1.],
        // w=[5 0 5 3 3 2 5 5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  78417.   24947.   50705.   97518.   -4669.  -14514.   80458. -100104.], 
        // Q{mac}=[76 24 49 95  0  0 78  0]

        sign=8'b01001000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000101, 8'b00000000, 8'b00000101, 8'b00000011, 8'b00000011, 8'b00000010, 8'b00000101, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 495: 
        // x=-128, 
        // s=[-1. -1. -1. -1. -1.  1.  1.  1.],
        // w=[1 2 4 4 4 4 6 7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  78545.   25203.   51217.   98030.   -4157.  -15026.   79690. -101000.], 
        // Q{mac}=[76 24 50 95  0  0 77  0]

        sign=8'b00000111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00000010, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000110, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 496: 
        // x=-128, 
        // s=[-1.  1.  1. -1. -1.  1.  1. -1.],
        // w=[ 9  3  8 10  7  4  0  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  79697.   24819.   50193.   99310.   -3261.  -15538.   79690. -100360.], 
        // Q{mac}=[77 24 49 96  0  0 77  0]

        sign=8'b01100110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001001, 8'b00000011, 8'b00001000, 8'b00001010, 8'b00000111, 8'b00000100, 8'b00000000, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 497: 
        // x=-128, 
        // s=[ 1. -1.  1. -1.  1. -1.  1. -1.],
        // w=[0 3 7 1 3 5 2 1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  79697.   25203.   49297.   99438.   -3645.  -14898.   79434. -100232.], 
        // Q{mac}=[77 24 48 97  0  0 77  0]

        sign=8'b10101010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000000, 8'b00000011, 8'b00000111, 8'b00000001, 8'b00000011, 8'b00000101, 8'b00000010, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 498: 
        // x=-128, 
        // s=[ 1.  1. -1. -1. -1.  1.  1. -1.],
        // w=[ 6  5  1  8 11  5  2  1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  78929.   24563.   49425.  100462.   -2237.  -15538.   79178. -100104.], 
        // Q{mac}=[77 23 48 98  0  0 77  0]

        sign=8'b11000110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000110, 8'b00000101, 8'b00000001, 8'b00001000, 8'b00001011, 8'b00000101, 8'b00000010, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 499: 
        // x=-128, 
        // s=[-1. -1.  1. -1. -1.  1.  1.  1.],
        // w=[3 5 8 1 3 2 0 1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  79313.   25203.   48401.  100590.   -1853.  -15794.   79178. -100232.], 
        // Q{mac}=[77 24 47 98  0  0 77  0]

        sign=8'b00100111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00000101, 8'b00001000, 8'b00000001, 8'b00000011, 8'b00000010, 8'b00000000, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 500: 
        // x=-128, 
        // s=[-1. -1. -1. -1. -1.  1.  1.  1.],
        // w=[ 5 10  2  9  7  3  4  6],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  79953.   26483.   48657.  101742.    -957.  -16178.   78666. -101000.], 
        // Q{mac}=[78 25 47 99  0  0 76  0]

        sign=8'b00000111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000101, 8'b00001010, 8'b00000010, 8'b00001001, 8'b00000111, 8'b00000011, 8'b00000100, 8'b00000110};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 501: 
        // x=-102, 
        // s=[ 1.  1. -1. -1.  1.  1.  1.  1.],
        // w=[ 0 16 26 19  4  9  6  8],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  79953.   24851.   51309.  103680.   -1365.  -17096.   78054. -101816.], 
        // Q{mac}=[ 78  24  50 101   0   0  76   0]

        sign=8'b11001111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000000, 8'b00010000, 8'b00011010, 8'b00010011, 8'b00000100, 8'b00001001, 8'b00000110, 8'b00001000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10011010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 502: 
        // x=-92, 
        // s=[ 1.  1. -1. -1. -1.  1.  1.  1.],
        // w=[12 12 21  6  8 11  5  4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  78849.   23747.   53241.  104232.    -629.  -18108.   77594. -102184.], 
        // Q{mac}=[ 77  23  51 101   0   0  75   0]

        sign=8'b11000111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001100, 8'b00001100, 8'b00010101, 8'b00000110, 8'b00001000, 8'b00001011, 8'b00000101, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10100100;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 503: 
        // x=-94, 
        // s=[ 1.  1. -1. -1.  1.  1.  1.  1.],
        // w=[11 27 23 18  5  6 10  7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  77815.   21209.   55403.  105924.   -1099.  -18672.   76654. -102842.], 
        // Q{mac}=[ 75  20  54 103   0   0  74   0]

        sign=8'b11001111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001011, 8'b00011011, 8'b00010111, 8'b00010010, 8'b00000101, 8'b00000110, 8'b00001010, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10100010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 504: 
        // x=-100, 
        // s=[ 1.  1. -1. -1. -1.  1. -1. -1.],
        // w=[ 9  0  6  9 13  7  1  4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  76915.   21209.   56003.  106824.     201.  -19372.   76754. -102442.], 
        // Q{mac}=[ 75  20  54 104   0   0  74   0]

        sign=8'b11000100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001001, 8'b00000000, 8'b00000110, 8'b00001001, 8'b00001101, 8'b00000111, 8'b00000001, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10011100;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 505: 
        // x=-121, 
        // s=[ 1. -1. -1. -1. -1. -1. -1.  1.],
        // w=[2 1 4 3 5 3 5 8],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  76673.   21330.   56487.  107187.     806.  -19009.   77359. -103410.], 
        // Q{mac}=[ 74  20  55 104   0   0  75   0]

        sign=8'b10000001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00000001, 8'b00000100, 8'b00000011, 8'b00000101, 8'b00000011, 8'b00000101, 8'b00001000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000111;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 506: 
        // x=-102, 
        // s=[ 1.  1. -1. -1.  1. -1.  1.  1.],
        // w=[ 0 17 20 16  8  1  8  0],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 7.66730e+04  1.95960e+04  5.85270e+04  1.08819e+05 -1.00000e+01   -1.89070e+04  7.65430e+04 -1.03410e+05], 
        // Q{mac}=[ 74  19  57 106   0   0  74   0]

        sign=8'b11001011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000000, 8'b00010001, 8'b00010100, 8'b00010000, 8'b00001000, 8'b00000001, 8'b00001000, 8'b00000000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10011010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 507: 
        // x=-123, 
        // s=[ 1.  1. -1. -1. -1.  1.  1.  1.],
        // w=[ 4  8 22  5  4  1  8  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  76181.   18612.   61233.  109434.     482.  -19030.   75559. -103656.], 
        // Q{mac}=[ 74  18  59 106   0   0  73   0]

        sign=8'b11000111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000100, 8'b00001000, 8'b00010110, 8'b00000101, 8'b00000100, 8'b00000001, 8'b00001000, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 508: 
        // x=-112, 
        // s=[ 1.  1. -1. -1.  1.  1.  1. -1.],
        // w=[ 2 17 11 16  1  1  1  4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  75957.   16708.   62465.  111226.     370.  -19142.   75447. -103208.], 
        // Q{mac}=[ 74  16  61 108   0   0  73   0]

        sign=8'b11001110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00010001, 8'b00001011, 8'b00010000, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10010000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 509: 
        // x=-23, 
        // s=[-1.  1. -1. -1.  1.  1.  1.  1.],
        // w=[ 2  4  7 15 14  3 12  6],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 7.60030e+04  1.66160e+04  6.26260e+04  1.11571e+05  4.80000e+01   -1.92110e+04  7.51710e+04 -1.03346e+05], 
        // Q{mac}=[ 74  16  61 108   0   0  73   0]

        sign=8'b01001111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00000100, 8'b00000111, 8'b00001111, 8'b00001110, 8'b00000011, 8'b00001100, 8'b00000110};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11101001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 510: 
        // x=-128, 
        // s=[ 1. -1.  1. -1. -1.  1. -1. -1.],
        // w=[3 1 4 6 9 6 2 4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  75619.   16744.   62114.  112339.    1200.  -19979.   75427. -102834.], 
        // Q{mac}=[ 73  16  60 109   1   0  73   0]

        sign=8'b10100100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00000001, 8'b00000100, 8'b00000110, 8'b00001001, 8'b00000110, 8'b00000010, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 511: 
        // x=-63, 
        // s=[-1. -1.  1.  1.  1. -1. -1.  1.],
        // w=[12 10 12  5 13  5  8  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  76375.   17374.   61358.  112024.     381.  -19664.   75931. -103023.], 
        // Q{mac}=[ 74  16  59 109   0   0  74   0]

        sign=8'b00111001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001100, 8'b00001010, 8'b00001100, 8'b00000101, 8'b00001101, 8'b00000101, 8'b00001000, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11000001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 512: 
        // x=-50, 
        // s=[ 1. -1.  1.  1. -1. -1.  1. -1.],
        // w=[ 3  4  0  3 25  4  3  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  76225.   17574.   61358.  111874.    1631.  -19464.   75781. -102773.], 
        // Q{mac}=[ 74  17  59 109   1   0  74   0]

        sign=8'b10110010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00000100, 8'b00000000, 8'b00000011, 8'b00011001, 8'b00000100, 8'b00000011, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11001110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 513: 
        // x=-115, 
        // s=[-1. -1. -1. -1.  1. -1.  1. -1.],
        // w=[ 8  1  3  5 15  4 11  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[ 7.71450e+04  1.76890e+04  6.17030e+04  1.12449e+05 -9.40000e+01   -1.90040e+04  7.45160e+04 -1.02428e+05], 
        // Q{mac}=[ 75  17  60 109   0   0  72   0]

        sign=8'b00001010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001000, 8'b00000001, 8'b00000011, 8'b00000101, 8'b00001111, 8'b00000100, 8'b00001011, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 514: 
        // x=-115, 
        // s=[-1. -1. -1. -1.  1. -1. -1.  1.],
        // w=[ 5  2 12  2 16  6  5  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  77720.   17919.   63083.  112679.   -1934.  -18314.   75091. -103003.], 
        // Q{mac}=[ 75  17  61 110   0   0  73   0]

        sign=8'b00001001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000101, 8'b00000010, 8'b00001100, 8'b00000010, 8'b00010000, 8'b00000110, 8'b00000101, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 515: 
        // x=-114, 
        // s=[ 1.  1. -1. -1.  1. -1. -1.  1.],
        // w=[ 1  5  4 10 20  6  1  8],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  77606.   17349.   63539.  113819.   -4214.  -17630.   75205. -103915.], 
        // Q{mac}=[ 75  16  62 111   0   0  73   0]

        sign=8'b11001001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00000101, 8'b00000100, 8'b00001010, 8'b00010100, 8'b00000110, 8'b00000001, 8'b00001000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 516: 
        // x=-119, 
        // s=[-1.  1. -1.  1.  1. -1.  1. -1.],
        // w=[ 1  5  1  3 19 12  8  4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  77725.   16754.   63658.  113462.   -6475.  -16202.   74253. -103439.], 
        // Q{mac}=[ 75  16  62 110   0   0  72   0]

        sign=8'b01011010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00000101, 8'b00000001, 8'b00000011, 8'b00010011, 8'b00001100, 8'b00001000, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 517: 
        // x=-116, 
        // s=[-1.  1.  1. -1. -1.  1.  1.  1.],
        // w=[ 7  8  1 10 10 13  8  4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  78537.   15826.   63542.  114622.   -5315.  -17710.   73325. -103903.], 
        // Q{mac}=[ 76  15  62 111   0   0  71   0]

        sign=8'b01100111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00001000, 8'b00000001, 8'b00001010, 8'b00001010, 8'b00001101, 8'b00001000, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001100;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 518: 
        // x=-115, 
        // s=[-1.  1. -1. -1.  1.  1.  1. -1.],
        // w=[9 5 1 9 7 5 3 2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  79572.   15251.   63657.  115657.   -6120.  -18285.   72980. -103673.], 
        // Q{mac}=[ 77  14  62 112   0   0  71   0]

        sign=8'b01001110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001001, 8'b00000101, 8'b00000001, 8'b00001001, 8'b00000111, 8'b00000101, 8'b00000011, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 519: 
        // x=-128, 
        // s=[ 1.  1. -1. -1. -1.  1.  1. -1.],
        // w=[0 1 8 7 4 2 3 3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  79572.   15123.   64681.  116553.   -5608.  -18541.   72596. -103289.], 
        // Q{mac}=[ 77  14  63 113   0   0  70   0]

        sign=8'b11000110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000000, 8'b00000001, 8'b00001000, 8'b00000111, 8'b00000100, 8'b00000010, 8'b00000011, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 520: 
        // x=-118, 
        // s=[-1.  1.  1. -1.  1.  1.  1.  1.],
        // w=[10  7  2  5  3  0  2  1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  80752.   14297.   64445.  117143.   -5962.  -18541.   72360. -103407.], 
        // Q{mac}=[ 78  13  62 114   0   0  70   0]

        sign=8'b01101111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001010, 8'b00000111, 8'b00000010, 8'b00000101, 8'b00000011, 8'b00000000, 8'b00000010, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 521: 
        // x=-63, 
        // s=[-1.  1. -1. -1.  1.  1.  1. -1.],
        // w=[17  6 10 13 12 13  6  6],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  81823.   13919.   65075.  117962.   -6718.  -19360.   71982. -103029.], 
        // Q{mac}=[ 79  13  63 115   0   0  70   0]

        sign=8'b01001110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00010001, 8'b00000110, 8'b00001010, 8'b00001101, 8'b00001100, 8'b00001101, 8'b00000110, 8'b00000110};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11000001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 522: 
        // x=-128, 
        // s=[ 1.  1. -1. -1. -1. -1. -1.  1.],
        // w=[3 5 3 8 8 8 2 5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  81439.   13279.   65459.  118986.   -5694.  -18336.   72238. -103669.], 
        // Q{mac}=[ 79  12  63 116   0   0  70   0]

        sign=8'b11000001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00000101, 8'b00000011, 8'b00001000, 8'b00001000, 8'b00001000, 8'b00000010, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 523: 
        // x=-6, 
        // s=[-1. -1.  1. -1. -1.  1.  1.  1.],
        // w=[12  1  9  9  5 12 14  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  81511.   13285.   65405.  119040.   -5664.  -18408.   72154. -103681.], 
        // Q{mac}=[ 79  12  63 116   0   0  70   0]

        sign=8'b00100111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001100, 8'b00000001, 8'b00001001, 8'b00001001, 8'b00000101, 8'b00001100, 8'b00001110, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11111010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 524: 
        // x=-33, 
        // s=[-1.  1. -1.  1.  1. -1.  1.  1.],
        // w=[15  1 14 10 50 40  0  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  82006.   13252.   65867.  118710.   -7314.  -17088.   72154. -103747.], 
        // Q{mac}=[ 80  12  64 115   0   0  70   0]

        sign=8'b01011011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001111, 8'b00000001, 8'b00001110, 8'b00001010, 8'b00110010, 8'b00101000, 8'b00000000, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11011111;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 525: 
        // x=-90, 
        // s=[-1.  1. -1.  1.  1. -1. -1. -1.],
        // w=[11  4  5  5 17 22  4  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  82996.   12892.   66317.  118260.   -8844.  -15108.   72514. -103297.], 
        // Q{mac}=[ 81  12  64 115   0   0  70   0]

        sign=8'b01011000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001011, 8'b00000100, 8'b00000101, 8'b00000101, 8'b00010001, 8'b00010110, 8'b00000100, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10100110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 526: 
        // x=-99, 
        // s=[-1.  1. -1. -1.  1.  1. -1. -1.],
        // w=[ 7  8  2 10  9  6  1  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  83689.   12100.   66515.  119250.   -9735.  -15702.   72613. -103000.], 
        // Q{mac}=[ 81  11  64 116   0   0  70   0]

        sign=8'b01001100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00001000, 8'b00000010, 8'b00001010, 8'b00001001, 8'b00000110, 8'b00000001, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10011101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 527: 
        // x=-103, 
        // s=[ 1. -1. -1. -1. -1. -1. -1. -1.],
        // w=[8 2 1 5 2 3 3 3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  82865.   12306.   66618.  119765.   -9529.  -15393.   72922. -102691.], 
        // Q{mac}=[ 80  12  65 116   0   0  71   0]

        sign=8'b10000000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001000, 8'b00000010, 8'b00000001, 8'b00000101, 8'b00000010, 8'b00000011, 8'b00000011, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10011001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 528: 
        // x=-98, 
        // s=[ 1.  1. -1. -1.  1. -1. -1.  1.],
        // w=[ 2  1 11 12  5  2  5  0],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  82669.   12208.   67696.  120941.  -10019.  -15197.   73412. -102691.], 
        // Q{mac}=[ 80  11  66 118   0   0  71   0]

        sign=8'b11001001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00000001, 8'b00001011, 8'b00001100, 8'b00000101, 8'b00000010, 8'b00000101, 8'b00000000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10011110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 529: 
        // x=-106, 
        // s=[-1.  1.  1. -1.  1. -1.  1.  1.],
        // w=[2 3 3 4 9 9 1 1],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  82881.   11890.   67378.  121365.  -10973.  -14243.   73306. -102797.], 
        // Q{mac}=[ 80  11  65 118   0   0  71   0]

        sign=8'b01101011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00000011, 8'b00000011, 8'b00000100, 8'b00001001, 8'b00001001, 8'b00000001, 8'b00000001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10010110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 530: 
        // x=-121, 
        // s=[ 1.  1. -1. -1.  1.  1.  1.  1.],
        // w=[ 5 10  9  9  4  3  2  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  82276.   10680.   68467.  122454.  -11457.  -14606.   73064. -103402.], 
        // Q{mac}=[ 80  10  66 119   0   0  71   0]

        sign=8'b11001111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000101, 8'b00001010, 8'b00001001, 8'b00001001, 8'b00000100, 8'b00000011, 8'b00000010, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000111;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 531: 
        // x=-99, 
        // s=[ 1. -1.  1. -1.  1.  1.  1. -1.],
        // w=[5 3 1 7 2 7 6 6],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  81781.   10977.   68368.  123147.  -11655.  -15299.   72470. -102808.], 
        // Q{mac}=[ 79  10  66 120   0   0  70   0]

        sign=8'b10101110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000101, 8'b00000011, 8'b00000001, 8'b00000111, 8'b00000010, 8'b00000111, 8'b00000110, 8'b00000110};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10011101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 532: 
        // x=-125, 
        // s=[-1. -1. -1. -1. -1. -1. -1.  1.],
        // w=[6 1 4 1 1 5 6 7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  82531.   11102.   68868.  123272.  -11530.  -14674.   73220. -103683.], 
        // Q{mac}=[ 80  10  67 120   0   0  71   0]

        sign=8'b00000001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000110, 8'b00000001, 8'b00000100, 8'b00000001, 8'b00000001, 8'b00000101, 8'b00000110, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000011;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 533: 
        // x=-103, 
        // s=[-1. -1. -1.  1. -1.  1.  1.  1.],
        // w=[ 3  9 10  0  5  4  0  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  82840.   12029.   69898.  123272.  -11015.  -15086.   73220. -104198.], 
        // Q{mac}=[ 80  11  68 120   0   0  71   0]

        sign=8'b00010111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00001001, 8'b00001010, 8'b00000000, 8'b00000101, 8'b00000100, 8'b00000000, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10011001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 534: 
        // x=22, 
        // s=[-1.  1. -1. -1.  1.  1.  1.  1.],
        // w=[ 9  3 11  7 19  7  9  3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  82642.   12095.   69656.  123118.  -10597.  -14932.   73418. -104132.], 
        // Q{mac}=[ 80  11  68 120   0   0  71   0]

        sign=8'b01001111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001001, 8'b00000011, 8'b00001011, 8'b00000111, 8'b00010011, 8'b00000111, 8'b00001001, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00010110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 535: 
        // x=-128, 
        // s=[-1. -1.  1.  1.  1. -1. -1. -1.],
        // w=[15  2  5  6  5  9 10  4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  84562.   12351.   69016.  122350.  -11237.  -13780.   74698. -103620.], 
        // Q{mac}=[ 82  12  67 119   0   0  72   0]

        sign=8'b00111000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001111, 8'b00000010, 8'b00000101, 8'b00000110, 8'b00000101, 8'b00001001, 8'b00001010, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 536: 
        // x=-7, 
        // s=[-1. -1.  1.  1.  1. -1. -1.  1.],
        // w=[10  2  3 28 33 34 16  0],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  84632.   12365.   68995.  122154.  -11468.  -13542.   74810. -103620.], 
        // Q{mac}=[ 82  12  67 119   0   0  73   0]

        sign=8'b00111001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001010, 8'b00000010, 8'b00000011, 8'b00011100, 8'b00100001, 8'b00100010, 8'b00010000, 8'b00000000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11111001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 537: 
        // x=-61, 
        // s=[ 1.  1.  1.  1.  1. -1. -1. -1.],
        // w=[ 9  5  6  5  0  4 17  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  84083.   12060.   68629.  121849.  -11468.  -13298.   75847. -103498.], 
        // Q{mac}=[ 82  11  67 118   0   0  74   0]

        sign=8'b11111000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001001, 8'b00000101, 8'b00000110, 8'b00000101, 8'b00000000, 8'b00000100, 8'b00010001, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11000011;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 538: 
        // x=-98, 
        // s=[ 1.  1. -1.  1.  1. -1. -1. -1.],
        // w=[14  0  1  2  0  1 23  6],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  82711.   12060.   68727.  121653.  -11468.  -13200.   78101. -102910.], 
        // Q{mac}=[ 80  11  67 118   0   0  76   0]

        sign=8'b11011000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001110, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000000, 8'b00000001, 8'b00010111, 8'b00000110};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10011110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 539: 
        // x=-114, 
        // s=[-1.  1. -1.  1. -1. -1.  1.  1.],
        // w=[5 0 3 3 4 3 4 9],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  83281.   12060.   69069.  121311.  -11012.  -12858.   77645. -103936.], 
        // Q{mac}=[ 81  11  67 118   0   0  75   0]

        sign=8'b01010011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000101, 8'b00000000, 8'b00000011, 8'b00000011, 8'b00000100, 8'b00000011, 8'b00000100, 8'b00001001};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 540: 
        // x=-117, 
        // s=[-1. -1.  1.  1. -1.  1. -1.  1.],
        // w=[10  8  3  0  5  2  7  0],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  84451.   12996.   68718.  121311.  -10427.  -13092.   78464. -103936.], 
        // Q{mac}=[ 82  12  67 118   0   0  76   0]

        sign=8'b00110101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001010, 8'b00001000, 8'b00000011, 8'b00000000, 8'b00000101, 8'b00000010, 8'b00000111, 8'b00000000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001011;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 541: 
        // x=-115, 
        // s=[-1. -1. -1. -1.  1. -1. -1.  1.],
        // w=[ 8  5  1  3  5 10  1  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  85371.   13571.   68833.  121656.  -11002.  -11942.   78579. -104511.], 
        // Q{mac}=[ 83  13  67 118   0   0  76   0]

        sign=8'b00001001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001000, 8'b00000101, 8'b00000001, 8'b00000011, 8'b00000101, 8'b00001010, 8'b00000001, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 542: 
        // x=-118, 
        // s=[ 1. -1. -1.  1. -1.  1.  1.  1.],
        // w=[ 1  3  4  0 10  4  2  0],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  85253.   13925.   69305.  121656.   -9822.  -12414.   78343. -104511.], 
        // Q{mac}=[ 83  13  67 118   0   0  76   0]

        sign=8'b10010111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000001, 8'b00000011, 8'b00000100, 8'b00000000, 8'b00001010, 8'b00000100, 8'b00000010, 8'b00000000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 543: 
        // x=-117, 
        // s=[ 1. -1. -1. -1. -1. -1. -1.  1.],
        // w=[0 4 5 6 4 5 3 0],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  85253.   14393.   69890.  122358.   -9354.  -11829.   78694. -104511.], 
        // Q{mac}=[ 83  14  68 119   0   0  76   0]

        sign=8'b10000001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000000, 8'b00000100, 8'b00000101, 8'b00000110, 8'b00000100, 8'b00000101, 8'b00000011, 8'b00000000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001011;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 544: 
        // x=-114, 
        // s=[-1.  1. -1.  1. -1. -1. -1.  1.],
        // w=[2 0 8 1 6 4 3 7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  85481.   14393.   70802.  122244.   -8670.  -11373.   79036. -105309.], 
        // Q{mac}=[ 83  14  69 119   0   0  77   0]

        sign=8'b01010001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00000000, 8'b00001000, 8'b00000001, 8'b00000110, 8'b00000100, 8'b00000011, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 545: 
        // x=-128, 
        // s=[-1.  1.  1. -1. -1. -1. -1. -1.],
        // w=[7 0 8 4 5 8 4 3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  86377.   14393.   69778.  122756.   -8030.  -10349.   79548. -104925.], 
        // Q{mac}=[ 84  14  68 119   0   0  77   0]

        sign=8'b01100000;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000111, 8'b00000000, 8'b00001000, 8'b00000100, 8'b00000101, 8'b00001000, 8'b00000100, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 546: 
        // x=-115, 
        // s=[ 1.  1. -1. -1.  1. -1.  1. -1.],
        // w=[0 5 7 4 3 9 0 3],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  86377.   13818.   70583.  123216.   -8375.   -9314.   79548. -104580.], 
        // Q{mac}=[ 84  13  68 120   0   0  77   0]

        sign=8'b11001010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000000, 8'b00000101, 8'b00000111, 8'b00000100, 8'b00000011, 8'b00001001, 8'b00000000, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10001101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 547: 
        // x=-31, 
        // s=[-1.  1. -1.  1.  1. -1.  1. -1.],
        // w=[14  2  5  7 22  5  2  4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  86811.   13756.   70738.  122999.   -9057.   -9159.   79486. -104456.], 
        // Q{mac}=[ 84  13  69 120   0   0  77   0]

        sign=8'b01011010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001110, 8'b00000010, 8'b00000101, 8'b00000111, 8'b00010110, 8'b00000101, 8'b00000010, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11100001;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 548: 
        // x=-128, 
        // s=[-1. -1. -1.  1.  1. -1.  1. -1.],
        // w=[8 6 7 5 2 7 3 4],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  87835.   14524.   71634.  122359.   -9313.   -8263.   79102. -103944.], 
        // Q{mac}=[ 85  14  69 119   0   0  77   0]

        sign=8'b00011010;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001000, 8'b00000110, 8'b00000111, 8'b00000101, 8'b00000010, 8'b00000111, 8'b00000011, 8'b00000100};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10000000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 549: 
        // x=8, 
        // s=[-1. -1.  1. -1.  1.  1.  1.  1.],
        // w=[18  8  3  6 11  0 10  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  87691.   14460.   71658.  122311.   -9225.   -8263.   79182. -103928.], 
        // Q{mac}=[ 85  14  69 119   0   0  77   0]

        sign=8'b00101111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00010010, 8'b00001000, 8'b00000011, 8'b00000110, 8'b00001011, 8'b00000000, 8'b00001010, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00001000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 550: 
        // x=-43, 
        // s=[-1. -1.  1.  1. -1.  1. -1.  1.],
        // w=[ 2 11 29 22 14  1 20  8],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  87777.   14933.   70411.  121365.   -8623.   -8306.   80042. -104272.], 
        // Q{mac}=[ 85  14  68 118   0   0  78   0]

        sign=8'b00110101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00001011, 8'b00011101, 8'b00010110, 8'b00001110, 8'b00000001, 8'b00010100, 8'b00001000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b11010101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 551: 
        // x=-91, 
        // s=[ 1. -1.  1.  1. -1.  1. -1. -1.],
        // w=[ 3 21 21 13  2  3  7  5],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  87504.   16844.   68500.  120182.   -8441.   -8579.   80679. -103817.], 
        // Q{mac}=[ 85  16  66 117   0   0  78   0]

        sign=8'b10110100;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000011, 8'b00010101, 8'b00010101, 8'b00001101, 8'b00000010, 8'b00000011, 8'b00000111, 8'b00000101};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10100101;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 552: 
        // x=20, 
        // s=[ 1. -1. -1.  1.  1. -1. -1.  1.],
        // w=[8 5 5 4 1 1 1 7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  87664.   16744.   68400.  120262.   -8421.   -8599.   80659. -103677.], 
        // Q{mac}=[ 85  16  66 117   0   0  78   0]

        sign=8'b10011001;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001000, 8'b00000101, 8'b00000101, 8'b00000100, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00010100;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 553: 
        // x=-106, 
        // s=[-1. -1. -1. -1.  1. -1.  1.  1.],
        // w=[13  2 10  4 16  4 22  0],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  89042.   16956.   69460.  120686.  -10117.   -8175.   78327. -103677.], 
        // Q{mac}=[ 86  16  67 117   0   0  76   0]

        sign=8'b00001011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001101, 8'b00000010, 8'b00001010, 8'b00000100, 8'b00010000, 8'b00000100, 8'b00010110, 8'b00000000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10010110;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 554: 
        // x=34, 
        // s=[-1. -1. -1.  1. -1. -1.  1.  1.],
        // w=[12  3 13  7  8  6  8  2],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  88634.   16854.   69018.  120924.  -10389.   -8379.   78599. -103609.], 
        // Q{mac}=[ 86  16  67 118   0   0  76   0]

        sign=8'b00010011;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00001100, 8'b00000011, 8'b00001101, 8'b00000111, 8'b00001000, 8'b00000110, 8'b00001000, 8'b00000010};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00100010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 555: 
        // x=-93, 
        // s=[ 1.  1. -1.  1. -1.  1. -1.  1.],
        // w=[34  2 65 38 19 16  8  8],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  85472.   16668.   75063.  117390.   -8622.   -9867.   79343. -104353.], 
        // Q{mac}=[ 83  16  73 114   0   0  77   0]

        sign=8'b11010101;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00100010, 8'b00000010, 8'b01000001, 8'b00100110, 8'b00010011, 8'b00010000, 8'b00001000, 8'b00001000};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b10100011;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 556: 
        // x=34, 
        // s=[-1. -1.  1. -1. -1.  1.  1. -1.],
        // w=[44 88 23  8 31 16 85  7],
        // bias=[0 0 0 0 0 0 0 0],
        // mac=[  83976.   13676.   75845.  117118.   -9676.   -9323.   82233. -104591.], 
        // Q{mac}=[ 82  13  74 114   0   0  80   0]

        sign=8'b00100110;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00101100, 8'b01011000, 8'b00010111, 8'b00001000, 8'b00011111, 8'b00010000, 8'b01010101, 8'b00000111};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
        din=8'b00100010;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------
        // Operation 557: 
        // x=-8, 
        // s=[-1. -1. -1.  1. -1.  1.  1.  1.],
        // w=[ 2 23  3 11 14 17 18  3],
        // bias=[ 118  127   44  127  127  127  127 -128],
        // mac=[  83992.   13860.   75869.  117030.   -9564.   -9459.   82089. -104615.], 
        //  

        sign=8'b00010111;
        {win0, win1, win2, win3, win4, win5, win6, win7}={8'b00000010, 8'b00010111, 8'b00000011, 8'b00001011, 8'b00001110, 8'b00010001, 8'b00010010, 8'b00000011};
        {bias0, bias1, bias2, bias3, bias4, bias5, bias6, bias7}={8'b01110110, 8'b01111111, 8'b00101100, 8'b01111111, 8'b01111111, 8'b01111111, 8'b01111111, 8'b10000000};
        din=8'b11111000;
        trig = 1;  // Activate trig
        #50 trig = 0;
        #100000;
        //wait for clk_period;
        //----------------------------------------------------------------



        // Finish simulation
        $finish;
    end

endmodule
